module CELL_TYPE_CONST #(parameter PARAM_WIDTH=1, parameter PARAM_INIT_VALUE=0) (output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT); assign PORT_ID_OUT = PARAM_INIT_VALUE;
endmodule

module CELL_TYPE_MUL #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT); assign PORT_ID_OUT = PORT_ID_IN0 * PORT_ID_IN1;
 endmodule

module CELL_TYPE_ADD #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT); assign PORT_ID_OUT = PORT_ID_IN0 + PORT_ID_IN1;
 endmodule

module CELL_TYPE_SUB #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT); assign PORT_ID_OUT = PORT_ID_IN0 - PORT_ID_IN1;
 endmodule

module CELL_TYPE_AND #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT); assign PORT_ID_OUT = PORT_ID_IN0 & PORT_ID_IN1;
 endmodule

module CELL_TYPE_OR #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT); assign PORT_ID_OUT = PORT_ID_IN0 | PORT_ID_IN1;
 endmodule

module CELL_TYPE_EQ #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [0 : 0] PORT_ID_OUT); assign PORT_ID_OUT = PORT_ID_IN0 == PORT_ID_IN1;
 endmodule

module CELL_TYPE_ULT #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [0 : 0] PORT_ID_OUT); assign PORT_ID_OUT = PORT_ID_IN0 < PORT_ID_IN1;
 endmodule

module CELL_TYPE_UGE #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [0 : 0] PORT_ID_OUT); assign PORT_ID_OUT = PORT_ID_IN0 >= PORT_ID_IN1;
endmodule // CELL_TYPE_UGE

module CELL_TYPE_REG #(parameter PARAM_CLK_POSEDGE=1, parameter PARAM_INIT_VALUE=0, parameter PARAM_WIDTH=1)(input PORT_ID_CLK, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT);

   reg [PARAM_WIDTH - 1 : 0] data;
   
   initial begin
      data = PARAM_INIT_VALUE;
   end

   wire true_clk;
   assign true_clk = PARAM_CLK_POSEDGE ? PORT_ID_CLK : ~PORT_ID_CLK;
   
   always @(posedge true_clk) begin
      data <= PORT_ID_IN;
   end

   assign PORT_ID_OUT = data;
   
endmodule

module CELL_TYPE_REG_ARST #(parameter PARAM_CLK_POSEDGE=1, parameter PARAM_ARST_POSEDGE=1, parameter PARAM_INIT_VALUE=0, parameter PARAM_WIDTH=1)(input PORT_ID_ARST, input PORT_ID_CLK, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT);
   assign PORT_ID_OUT = 0;
   
endmodule // CELL_TYPE_REG_ARST

module CELL_TYPE_MEM #(parameter PARAM_HAS_INIT=0, parameter PARAM_MEM_DEPTH=0, parameter PARAM_MEM_WIDTH=0)(input PORT_ID_ARST, input PORT_ID_CLK, input PORT_ID_WEN, input [$clog2(PARAM_MEM_DEPTH) - 1 : 0] PORT_ID_RADDR, input [$clog2(PARAM_MEM_DEPTH) - 1 : 0] PORT_ID_WADDR, input [PARAM_MEM_WIDTH - 1 : 0] PORT_ID_WDATA, output [PARAM_MEM_WIDTH - 1 : 0] PORT_ID_RDATA);
   
   assign PORT_ID_RDATA = 0;
   
endmodule

module CELL_TYPE_MUX #(parameter PARAM_WIDTH=1) (input PORT_ID_SEL, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT);
   assign PORT_ID_OUT = PORT_ID_SEL ? PORT_ID_IN1 : PORT_ID_IN0;
 endmodule

module CELL_TYPE_NOT #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT); assign PORT_ID_OUT = ~PORT_ID_IN;
 endmodule

module CELL_TYPE_ORR #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT); assign PORT_ID_OUT = |PORT_ID_IN;
 endmodule

module CELL_TYPE_PORT #(parameter PARAM_PORT_TYPE=0, parameter PARAM_OUT_WIDTH=1) (input [PARAM_OUT_WIDTH - 1 : 0] PORT_ID_IN, output [PARAM_OUT_WIDTH - 1 : 0] PORT_ID_OUT); assign PORT_ID_OUT = PORT_ID_IN;
 endmodule

module CELL_TYPE_ZEXT #(parameter PARAM_IN_WIDTH=1, parameter PARAM_OUT_WIDTH=1) (input [PARAM_IN_WIDTH - 1 : 0] PORT_ID_IN, output [PARAM_OUT_WIDTH - 1 : 0] PORT_ID_OUT); assign PORT_ID_OUT = {{(PARAM_OUT_WIDTH - PARAM_IN_WIDTH){1'b0}}, PORT_ID_IN};
 endmodule


module top(	output [0 : 0] aux_div_pad,
	input [0 : 0] clk_ext_in,
	input [0 : 0] clk_in,
	input [31 : 0] config_addr_in,
	input [31 : 0] config_data_in,
	input [0 : 0] ext_cki,
	input [0 : 0] ext_cki_jm,
	input [0 : 0] ext_ckib,
	input [0 : 0] ext_ckib_jm,
	input [0 : 0] ext_frefn,
	input [0 : 0] ext_frefn_jm,
	input [0 : 0] ext_frefp,
	input [0 : 0] ext_frefp_jm,
	output [0 : 0] ffeed_pad,
	output [0 : 0] fout_div_pad,
	output [0 : 0] fref_off_pad,
	output [0 : 0] frefn_out_jm,
	output [0 : 0] frefp_out_jm,
	output [12 : 0] lf_out,
	output [3 : 0] mdllout_pad,
	input [0 : 0] pad_S0_T0_in,
	output [0 : 0] pad_S0_T0_out,
	input [0 : 0] pad_S0_T10_in,
	output [0 : 0] pad_S0_T10_out,
	input [0 : 0] pad_S0_T11_in,
	output [0 : 0] pad_S0_T11_out,
	input [0 : 0] pad_S0_T12_in,
	output [0 : 0] pad_S0_T12_out,
	input [0 : 0] pad_S0_T13_in,
	output [0 : 0] pad_S0_T13_out,
	input [0 : 0] pad_S0_T14_in,
	output [0 : 0] pad_S0_T14_out,
	input [0 : 0] pad_S0_T15_in,
	output [0 : 0] pad_S0_T15_out,
	input [0 : 0] pad_S0_T1_in,
	output [0 : 0] pad_S0_T1_out,
	input [0 : 0] pad_S0_T2_in,
	output [0 : 0] pad_S0_T2_out,
	input [0 : 0] pad_S0_T3_in,
	output [0 : 0] pad_S0_T3_out,
	input [0 : 0] pad_S0_T4_in,
	output [0 : 0] pad_S0_T4_out,
	input [0 : 0] pad_S0_T5_in,
	output [0 : 0] pad_S0_T5_out,
	input [0 : 0] pad_S0_T6_in,
	output [0 : 0] pad_S0_T6_out,
	input [0 : 0] pad_S0_T7_in,
	output [0 : 0] pad_S0_T7_out,
	input [0 : 0] pad_S0_T8_in,
	output [0 : 0] pad_S0_T8_out,
	input [0 : 0] pad_S0_T9_in,
	output [0 : 0] pad_S0_T9_out,
	input [0 : 0] pad_S1_T0_in,
	output [0 : 0] pad_S1_T0_out,
	input [0 : 0] pad_S1_T10_in,
	output [0 : 0] pad_S1_T10_out,
	input [0 : 0] pad_S1_T11_in,
	output [0 : 0] pad_S1_T11_out,
	input [0 : 0] pad_S1_T12_in,
	output [0 : 0] pad_S1_T12_out,
	input [0 : 0] pad_S1_T13_in,
	output [0 : 0] pad_S1_T13_out,
	input [0 : 0] pad_S1_T14_in,
	output [0 : 0] pad_S1_T14_out,
	input [0 : 0] pad_S1_T15_in,
	output [0 : 0] pad_S1_T15_out,
	input [0 : 0] pad_S1_T1_in,
	output [0 : 0] pad_S1_T1_out,
	input [0 : 0] pad_S1_T2_in,
	output [0 : 0] pad_S1_T2_out,
	input [0 : 0] pad_S1_T3_in,
	output [0 : 0] pad_S1_T3_out,
	input [0 : 0] pad_S1_T4_in,
	output [0 : 0] pad_S1_T4_out,
	input [0 : 0] pad_S1_T5_in,
	output [0 : 0] pad_S1_T5_out,
	input [0 : 0] pad_S1_T6_in,
	output [0 : 0] pad_S1_T6_out,
	input [0 : 0] pad_S1_T7_in,
	output [0 : 0] pad_S1_T7_out,
	input [0 : 0] pad_S1_T8_in,
	output [0 : 0] pad_S1_T8_out,
	input [0 : 0] pad_S1_T9_in,
	output [0 : 0] pad_S1_T9_out,
	input [0 : 0] pad_S2_T0_in,
	output [0 : 0] pad_S2_T0_out,
	input [0 : 0] pad_S2_T10_in,
	output [0 : 0] pad_S2_T10_out,
	input [0 : 0] pad_S2_T11_in,
	output [0 : 0] pad_S2_T11_out,
	input [0 : 0] pad_S2_T12_in,
	output [0 : 0] pad_S2_T12_out,
	input [0 : 0] pad_S2_T13_in,
	output [0 : 0] pad_S2_T13_out,
	input [0 : 0] pad_S2_T14_in,
	output [0 : 0] pad_S2_T14_out,
	input [0 : 0] pad_S2_T15_in,
	output [0 : 0] pad_S2_T15_out,
	input [0 : 0] pad_S2_T1_in,
	output [0 : 0] pad_S2_T1_out,
	input [0 : 0] pad_S2_T2_in,
	output [0 : 0] pad_S2_T2_out,
	input [0 : 0] pad_S2_T3_in,
	output [0 : 0] pad_S2_T3_out,
	input [0 : 0] pad_S2_T4_in,
	output [0 : 0] pad_S2_T4_out,
	input [0 : 0] pad_S2_T5_in,
	output [0 : 0] pad_S2_T5_out,
	input [0 : 0] pad_S2_T6_in,
	output [0 : 0] pad_S2_T6_out,
	input [0 : 0] pad_S2_T7_in,
	output [0 : 0] pad_S2_T7_out,
	input [0 : 0] pad_S2_T8_in,
	output [0 : 0] pad_S2_T8_out,
	input [0 : 0] pad_S2_T9_in,
	output [0 : 0] pad_S2_T9_out,
	input [0 : 0] pad_S3_T0_in,
	output [0 : 0] pad_S3_T0_out,
	input [0 : 0] pad_S3_T10_in,
	output [0 : 0] pad_S3_T10_out,
	input [0 : 0] pad_S3_T11_in,
	output [0 : 0] pad_S3_T11_out,
	input [0 : 0] pad_S3_T12_in,
	output [0 : 0] pad_S3_T12_out,
	input [0 : 0] pad_S3_T13_in,
	output [0 : 0] pad_S3_T13_out,
	input [0 : 0] pad_S3_T14_in,
	output [0 : 0] pad_S3_T14_out,
	input [0 : 0] pad_S3_T15_in,
	output [0 : 0] pad_S3_T15_out,
	input [0 : 0] pad_S3_T1_in,
	output [0 : 0] pad_S3_T1_out,
	input [0 : 0] pad_S3_T2_in,
	output [0 : 0] pad_S3_T2_out,
	input [0 : 0] pad_S3_T3_in,
	output [0 : 0] pad_S3_T3_out,
	input [0 : 0] pad_S3_T4_in,
	output [0 : 0] pad_S3_T4_out,
	input [0 : 0] pad_S3_T5_in,
	output [0 : 0] pad_S3_T5_out,
	input [0 : 0] pad_S3_T6_in,
	output [0 : 0] pad_S3_T6_out,
	input [0 : 0] pad_S3_T7_in,
	output [0 : 0] pad_S3_T7_out,
	input [0 : 0] pad_S3_T8_in,
	output [0 : 0] pad_S3_T8_out,
	input [0 : 0] pad_S3_T9_in,
	output [0 : 0] pad_S3_T9_out,
	input [0 : 0] reset_in,
	input [0 : 0] tck,
	input [0 : 0] tdi,
	output [0 : 0] tdo,
	input [0 : 0] tms,
	input [0 : 0] trst_n);

	wire [0 : 0] fresh_wire_0;
	wire [0 : 0] fresh_wire_1;
	wire [0 : 0] fresh_wire_2;
	wire [31 : 0] fresh_wire_3;
	wire [31 : 0] fresh_wire_4;
	wire [0 : 0] fresh_wire_5;
	wire [0 : 0] fresh_wire_6;
	wire [0 : 0] fresh_wire_7;
	wire [0 : 0] fresh_wire_8;
	wire [0 : 0] fresh_wire_9;
	wire [0 : 0] fresh_wire_10;
	wire [0 : 0] fresh_wire_11;
	wire [0 : 0] fresh_wire_12;
	wire [0 : 0] fresh_wire_13;
	wire [0 : 0] fresh_wire_14;
	wire [0 : 0] fresh_wire_15;
	wire [0 : 0] fresh_wire_16;
	wire [0 : 0] fresh_wire_17;
	wire [12 : 0] fresh_wire_18;
	wire [3 : 0] fresh_wire_19;
	wire [0 : 0] fresh_wire_20;
	wire [0 : 0] fresh_wire_21;
	wire [0 : 0] fresh_wire_22;
	wire [0 : 0] fresh_wire_23;
	wire [0 : 0] fresh_wire_24;
	wire [0 : 0] fresh_wire_25;
	wire [0 : 0] fresh_wire_26;
	wire [0 : 0] fresh_wire_27;
	wire [0 : 0] fresh_wire_28;
	wire [0 : 0] fresh_wire_29;
	wire [0 : 0] fresh_wire_30;
	wire [0 : 0] fresh_wire_31;
	wire [0 : 0] fresh_wire_32;
	wire [0 : 0] fresh_wire_33;
	wire [0 : 0] fresh_wire_34;
	wire [0 : 0] fresh_wire_35;
	wire [0 : 0] fresh_wire_36;
	wire [0 : 0] fresh_wire_37;
	wire [0 : 0] fresh_wire_38;
	wire [0 : 0] fresh_wire_39;
	wire [0 : 0] fresh_wire_40;
	wire [0 : 0] fresh_wire_41;
	wire [0 : 0] fresh_wire_42;
	wire [0 : 0] fresh_wire_43;
	wire [0 : 0] fresh_wire_44;
	wire [0 : 0] fresh_wire_45;
	wire [0 : 0] fresh_wire_46;
	wire [0 : 0] fresh_wire_47;
	wire [0 : 0] fresh_wire_48;
	wire [0 : 0] fresh_wire_49;
	wire [0 : 0] fresh_wire_50;
	wire [0 : 0] fresh_wire_51;
	wire [0 : 0] fresh_wire_52;
	wire [0 : 0] fresh_wire_53;
	wire [0 : 0] fresh_wire_54;
	wire [0 : 0] fresh_wire_55;
	wire [0 : 0] fresh_wire_56;
	wire [0 : 0] fresh_wire_57;
	wire [0 : 0] fresh_wire_58;
	wire [0 : 0] fresh_wire_59;
	wire [0 : 0] fresh_wire_60;
	wire [0 : 0] fresh_wire_61;
	wire [0 : 0] fresh_wire_62;
	wire [0 : 0] fresh_wire_63;
	wire [0 : 0] fresh_wire_64;
	wire [0 : 0] fresh_wire_65;
	wire [0 : 0] fresh_wire_66;
	wire [0 : 0] fresh_wire_67;
	wire [0 : 0] fresh_wire_68;
	wire [0 : 0] fresh_wire_69;
	wire [0 : 0] fresh_wire_70;
	wire [0 : 0] fresh_wire_71;
	wire [0 : 0] fresh_wire_72;
	wire [0 : 0] fresh_wire_73;
	wire [0 : 0] fresh_wire_74;
	wire [0 : 0] fresh_wire_75;
	wire [0 : 0] fresh_wire_76;
	wire [0 : 0] fresh_wire_77;
	wire [0 : 0] fresh_wire_78;
	wire [0 : 0] fresh_wire_79;
	wire [0 : 0] fresh_wire_80;
	wire [0 : 0] fresh_wire_81;
	wire [0 : 0] fresh_wire_82;
	wire [0 : 0] fresh_wire_83;
	wire [0 : 0] fresh_wire_84;
	wire [0 : 0] fresh_wire_85;
	wire [0 : 0] fresh_wire_86;
	wire [0 : 0] fresh_wire_87;
	wire [0 : 0] fresh_wire_88;
	wire [0 : 0] fresh_wire_89;
	wire [0 : 0] fresh_wire_90;
	wire [0 : 0] fresh_wire_91;
	wire [0 : 0] fresh_wire_92;
	wire [0 : 0] fresh_wire_93;
	wire [0 : 0] fresh_wire_94;
	wire [0 : 0] fresh_wire_95;
	wire [0 : 0] fresh_wire_96;
	wire [0 : 0] fresh_wire_97;
	wire [0 : 0] fresh_wire_98;
	wire [0 : 0] fresh_wire_99;
	wire [0 : 0] fresh_wire_100;
	wire [0 : 0] fresh_wire_101;
	wire [0 : 0] fresh_wire_102;
	wire [0 : 0] fresh_wire_103;
	wire [0 : 0] fresh_wire_104;
	wire [0 : 0] fresh_wire_105;
	wire [0 : 0] fresh_wire_106;
	wire [0 : 0] fresh_wire_107;
	wire [0 : 0] fresh_wire_108;
	wire [0 : 0] fresh_wire_109;
	wire [0 : 0] fresh_wire_110;
	wire [0 : 0] fresh_wire_111;
	wire [0 : 0] fresh_wire_112;
	wire [0 : 0] fresh_wire_113;
	wire [0 : 0] fresh_wire_114;
	wire [0 : 0] fresh_wire_115;
	wire [0 : 0] fresh_wire_116;
	wire [0 : 0] fresh_wire_117;
	wire [0 : 0] fresh_wire_118;
	wire [0 : 0] fresh_wire_119;
	wire [0 : 0] fresh_wire_120;
	wire [0 : 0] fresh_wire_121;
	wire [0 : 0] fresh_wire_122;
	wire [0 : 0] fresh_wire_123;
	wire [0 : 0] fresh_wire_124;
	wire [0 : 0] fresh_wire_125;
	wire [0 : 0] fresh_wire_126;
	wire [0 : 0] fresh_wire_127;
	wire [0 : 0] fresh_wire_128;
	wire [0 : 0] fresh_wire_129;
	wire [0 : 0] fresh_wire_130;
	wire [0 : 0] fresh_wire_131;
	wire [0 : 0] fresh_wire_132;
	wire [0 : 0] fresh_wire_133;
	wire [0 : 0] fresh_wire_134;
	wire [0 : 0] fresh_wire_135;
	wire [0 : 0] fresh_wire_136;
	wire [0 : 0] fresh_wire_137;
	wire [0 : 0] fresh_wire_138;
	wire [0 : 0] fresh_wire_139;
	wire [0 : 0] fresh_wire_140;
	wire [0 : 0] fresh_wire_141;
	wire [0 : 0] fresh_wire_142;
	wire [0 : 0] fresh_wire_143;
	wire [0 : 0] fresh_wire_144;
	wire [0 : 0] fresh_wire_145;
	wire [0 : 0] fresh_wire_146;
	wire [0 : 0] fresh_wire_147;
	wire [0 : 0] fresh_wire_148;
	wire [0 : 0] fresh_wire_149;
	wire [0 : 0] fresh_wire_150;
	wire [0 : 0] fresh_wire_151;
	wire [0 : 0] fresh_wire_152;
	wire [0 : 0] fresh_wire_153;
	wire [12 : 0] fresh_wire_154;
	wire [0 : 0] fresh_wire_155;
	wire [0 : 0] fresh_wire_156;
	wire [0 : 0] fresh_wire_157;
	wire [0 : 0] fresh_wire_158;
	wire [0 : 0] fresh_wire_159;
	wire [0 : 0] fresh_wire_160;
	wire [0 : 0] fresh_wire_161;
	wire [0 : 0] fresh_wire_162;
	wire [0 : 0] fresh_wire_163;
	wire [15 : 0] fresh_wire_164;
	wire [15 : 0] fresh_wire_165;
	wire [15 : 0] fresh_wire_166;
	wire [1 : 0] fresh_wire_167;
	wire [15 : 0] fresh_wire_168;
	wire [15 : 0] fresh_wire_169;
	wire [15 : 0] fresh_wire_170;
	wire [15 : 0] fresh_wire_171;
	wire [15 : 0] fresh_wire_172;
	wire [31 : 0] fresh_wire_173;
	wire [31 : 0] fresh_wire_174;
	wire [31 : 0] fresh_wire_175;
	wire [31 : 0] fresh_wire_176;
	wire [15 : 0] fresh_wire_177;
	wire [31 : 0] fresh_wire_178;
	wire [31 : 0] fresh_wire_179;
	wire [31 : 0] fresh_wire_180;
	wire [31 : 0] fresh_wire_181;
	wire [15 : 0] fresh_wire_182;
	wire [31 : 0] fresh_wire_183;
	wire [31 : 0] fresh_wire_184;
	wire [31 : 0] fresh_wire_185;
	wire [31 : 0] fresh_wire_186;
	wire [15 : 0] fresh_wire_187;
	wire [15 : 0] fresh_wire_188;
	wire [15 : 0] fresh_wire_189;
	wire [15 : 0] fresh_wire_190;
	wire [15 : 0] fresh_wire_191;
	wire [15 : 0] fresh_wire_192;
	wire [15 : 0] fresh_wire_193;
	wire [15 : 0] fresh_wire_194;
	wire [15 : 0] fresh_wire_195;
	wire [15 : 0] fresh_wire_196;
	wire [15 : 0] fresh_wire_197;
	wire [15 : 0] fresh_wire_198;
	wire [0 : 0] fresh_wire_199;
	wire [0 : 0] fresh_wire_200;
	wire [0 : 0] fresh_wire_201;
	wire [1 : 0] fresh_wire_202;
	wire [1 : 0] fresh_wire_203;
	wire [0 : 0] fresh_wire_204;
	wire [1 : 0] fresh_wire_205;
	wire [1 : 0] fresh_wire_206;
	wire [0 : 0] fresh_wire_207;
	wire [1 : 0] fresh_wire_208;
	wire [1 : 0] fresh_wire_209;
	wire [0 : 0] fresh_wire_210;
	wire [15 : 0] fresh_wire_211;
	wire [15 : 0] fresh_wire_212;
	wire [0 : 0] fresh_wire_213;
	wire [0 : 0] fresh_wire_214;
	wire [0 : 0] fresh_wire_215;
	wire [0 : 0] fresh_wire_216;
	wire [0 : 0] fresh_wire_217;
	wire [0 : 0] fresh_wire_218;
	wire [0 : 0] fresh_wire_219;
	wire [0 : 0] fresh_wire_220;
	wire [0 : 0] fresh_wire_221;
	wire [0 : 0] fresh_wire_222;
	wire [0 : 0] fresh_wire_223;
	wire [0 : 0] fresh_wire_224;
	wire [0 : 0] fresh_wire_225;
	wire [1 : 0] fresh_wire_226;
	wire [1 : 0] fresh_wire_227;
	wire [0 : 0] fresh_wire_228;
	wire [0 : 0] fresh_wire_229;
	wire [0 : 0] fresh_wire_230;
	wire [0 : 0] fresh_wire_231;
	wire [0 : 0] fresh_wire_232;
	wire [0 : 0] fresh_wire_233;
	wire [0 : 0] fresh_wire_234;
	wire [1 : 0] fresh_wire_235;
	wire [1 : 0] fresh_wire_236;
	wire [0 : 0] fresh_wire_237;
	wire [0 : 0] fresh_wire_238;
	wire [0 : 0] fresh_wire_239;
	wire [0 : 0] fresh_wire_240;
	wire [0 : 0] fresh_wire_241;
	wire [0 : 0] fresh_wire_242;
	wire [0 : 0] fresh_wire_243;
	wire [1 : 0] fresh_wire_244;
	wire [1 : 0] fresh_wire_245;
	wire [0 : 0] fresh_wire_246;
	wire [1 : 0] fresh_wire_247;
	wire [1 : 0] fresh_wire_248;
	wire [0 : 0] fresh_wire_249;
	wire [15 : 0] fresh_wire_250;
	wire [15 : 0] fresh_wire_251;
	wire [0 : 0] fresh_wire_252;
	wire [0 : 0] fresh_wire_253;
	wire [0 : 0] fresh_wire_254;
	wire [0 : 0] fresh_wire_255;
	wire [0 : 0] fresh_wire_256;
	wire [0 : 0] fresh_wire_257;
	wire [0 : 0] fresh_wire_258;
	wire [15 : 0] fresh_wire_259;
	wire [15 : 0] fresh_wire_260;
	wire [0 : 0] fresh_wire_261;
	wire [15 : 0] fresh_wire_262;
	wire [15 : 0] fresh_wire_263;
	wire [0 : 0] fresh_wire_264;
	wire [15 : 0] fresh_wire_265;
	wire [15 : 0] fresh_wire_266;
	wire [0 : 0] fresh_wire_267;
	wire [0 : 0] fresh_wire_268;
	wire [0 : 0] fresh_wire_269;
	wire [0 : 0] fresh_wire_270;
	wire [0 : 0] fresh_wire_271;
	wire [0 : 0] fresh_wire_272;
	wire [0 : 0] fresh_wire_273;
	wire [0 : 0] fresh_wire_274;
	wire [0 : 0] fresh_wire_275;
	wire [0 : 0] fresh_wire_276;
	wire [0 : 0] fresh_wire_277;
	wire [0 : 0] fresh_wire_278;
	wire [0 : 0] fresh_wire_279;
	wire [0 : 0] fresh_wire_280;
	wire [0 : 0] fresh_wire_281;
	wire [0 : 0] fresh_wire_282;
	wire [0 : 0] fresh_wire_283;
	wire [0 : 0] fresh_wire_284;
	wire [0 : 0] fresh_wire_285;
	wire [0 : 0] fresh_wire_286;
	wire [0 : 0] fresh_wire_287;
	wire [0 : 0] fresh_wire_288;
	wire [0 : 0] fresh_wire_289;
	wire [0 : 0] fresh_wire_290;
	wire [0 : 0] fresh_wire_291;
	wire [0 : 0] fresh_wire_292;
	wire [0 : 0] fresh_wire_293;
	wire [0 : 0] fresh_wire_294;
	wire [0 : 0] fresh_wire_295;
	wire [0 : 0] fresh_wire_296;
	wire [0 : 0] fresh_wire_297;
	wire [0 : 0] fresh_wire_298;
	wire [0 : 0] fresh_wire_299;
	wire [0 : 0] fresh_wire_300;
	wire [0 : 0] fresh_wire_301;
	wire [0 : 0] fresh_wire_302;
	wire [0 : 0] fresh_wire_303;
	wire [0 : 0] fresh_wire_304;
	wire [0 : 0] fresh_wire_305;
	wire [0 : 0] fresh_wire_306;
	wire [0 : 0] fresh_wire_307;
	wire [0 : 0] fresh_wire_308;
	wire [0 : 0] fresh_wire_309;
	wire [0 : 0] fresh_wire_310;
	wire [0 : 0] fresh_wire_311;
	wire [0 : 0] fresh_wire_312;
	wire [0 : 0] fresh_wire_313;
	wire [0 : 0] fresh_wire_314;
	wire [0 : 0] fresh_wire_315;
	wire [0 : 0] fresh_wire_316;
	wire [0 : 0] fresh_wire_317;
	wire [0 : 0] fresh_wire_318;
	wire [0 : 0] fresh_wire_319;
	wire [0 : 0] fresh_wire_320;
	wire [0 : 0] fresh_wire_321;
	wire [0 : 0] fresh_wire_322;
	wire [0 : 0] fresh_wire_323;
	wire [0 : 0] fresh_wire_324;
	wire [0 : 0] fresh_wire_325;
	wire [0 : 0] fresh_wire_326;
	wire [0 : 0] fresh_wire_327;
	wire [0 : 0] fresh_wire_328;
	wire [0 : 0] fresh_wire_329;
	wire [0 : 0] fresh_wire_330;
	wire [0 : 0] fresh_wire_331;
	wire [0 : 0] fresh_wire_332;
	wire [0 : 0] fresh_wire_333;
	wire [0 : 0] fresh_wire_334;
	wire [0 : 0] fresh_wire_335;
	wire [0 : 0] fresh_wire_336;
	wire [0 : 0] fresh_wire_337;
	wire [0 : 0] fresh_wire_338;
	wire [0 : 0] fresh_wire_339;
	wire [0 : 0] fresh_wire_340;
	wire [0 : 0] fresh_wire_341;
	wire [0 : 0] fresh_wire_342;
	wire [0 : 0] fresh_wire_343;
	wire [0 : 0] fresh_wire_344;
	wire [0 : 0] fresh_wire_345;
	wire [0 : 0] fresh_wire_346;
	wire [0 : 0] fresh_wire_347;
	wire [0 : 0] fresh_wire_348;
	wire [0 : 0] fresh_wire_349;
	wire [0 : 0] fresh_wire_350;
	wire [0 : 0] fresh_wire_351;
	wire [0 : 0] fresh_wire_352;
	wire [0 : 0] fresh_wire_353;
	wire [0 : 0] fresh_wire_354;
	wire [0 : 0] fresh_wire_355;
	wire [0 : 0] fresh_wire_356;
	wire [0 : 0] fresh_wire_357;
	wire [0 : 0] fresh_wire_358;
	wire [0 : 0] fresh_wire_359;
	wire [0 : 0] fresh_wire_360;
	wire [15 : 0] fresh_wire_361;
	wire [15 : 0] fresh_wire_362;
	wire [0 : 0] fresh_wire_363;
	wire [15 : 0] fresh_wire_364;
	wire [15 : 0] fresh_wire_365;
	wire [0 : 0] fresh_wire_366;
	wire [0 : 0] fresh_wire_367;
	wire [0 : 0] fresh_wire_368;
	wire [0 : 0] fresh_wire_369;
	wire [0 : 0] fresh_wire_370;
	wire [0 : 0] fresh_wire_371;
	wire [1 : 0] fresh_wire_372;
	wire [1 : 0] fresh_wire_373;
	wire [0 : 0] fresh_wire_374;
	wire [1 : 0] fresh_wire_375;
	wire [1 : 0] fresh_wire_376;
	wire [0 : 0] fresh_wire_377;
	wire [15 : 0] fresh_wire_378;
	wire [15 : 0] fresh_wire_379;
	wire [0 : 0] fresh_wire_380;
	wire [0 : 0] fresh_wire_381;
	wire [0 : 0] fresh_wire_382;
	wire [0 : 0] fresh_wire_383;
	wire [0 : 0] fresh_wire_384;
	wire [0 : 0] fresh_wire_385;
	wire [0 : 0] fresh_wire_386;
	wire [0 : 0] fresh_wire_387;
	wire [0 : 0] fresh_wire_388;
	wire [0 : 0] fresh_wire_389;
	wire [0 : 0] fresh_wire_390;
	wire [0 : 0] fresh_wire_391;
	wire [0 : 0] fresh_wire_392;
	wire [0 : 0] fresh_wire_393;
	wire [0 : 0] fresh_wire_394;
	wire [0 : 0] fresh_wire_395;
	wire [0 : 0] fresh_wire_396;
	wire [0 : 0] fresh_wire_397;
	wire [0 : 0] fresh_wire_398;
	wire [0 : 0] fresh_wire_399;
	wire [0 : 0] fresh_wire_400;
	wire [1 : 0] fresh_wire_401;
	wire [1 : 0] fresh_wire_402;
	wire [0 : 0] fresh_wire_403;
	wire [0 : 0] fresh_wire_404;
	wire [15 : 0] fresh_wire_405;
	wire [15 : 0] fresh_wire_406;
	wire [0 : 0] fresh_wire_407;
	wire [0 : 0] fresh_wire_408;
	wire [15 : 0] fresh_wire_409;
	wire [15 : 0] fresh_wire_410;
	wire [0 : 0] fresh_wire_411;
	wire [0 : 0] fresh_wire_412;
	wire [15 : 0] fresh_wire_413;
	wire [15 : 0] fresh_wire_414;
	wire [0 : 0] fresh_wire_415;
	wire [0 : 0] fresh_wire_416;
	wire [15 : 0] fresh_wire_417;
	wire [15 : 0] fresh_wire_418;
	wire [0 : 0] fresh_wire_419;
	wire [0 : 0] fresh_wire_420;
	wire [0 : 0] fresh_wire_421;
	wire [0 : 0] fresh_wire_422;
	wire [0 : 0] fresh_wire_423;
	wire [0 : 0] fresh_wire_424;
	wire [0 : 0] fresh_wire_425;
	wire [0 : 0] fresh_wire_426;
	wire [0 : 0] fresh_wire_427;
	wire [0 : 0] fresh_wire_428;
	wire [0 : 0] fresh_wire_429;
	wire [0 : 0] fresh_wire_430;
	wire [0 : 0] fresh_wire_431;
	wire [0 : 0] fresh_wire_432;
	wire [15 : 0] fresh_wire_433;
	wire [15 : 0] fresh_wire_434;
	wire [15 : 0] fresh_wire_435;
	wire [0 : 0] fresh_wire_436;
	wire [0 : 0] fresh_wire_437;
	wire [0 : 0] fresh_wire_438;
	wire [0 : 0] fresh_wire_439;
	wire [0 : 0] fresh_wire_440;
	wire [0 : 0] fresh_wire_441;
	wire [0 : 0] fresh_wire_442;
	wire [0 : 0] fresh_wire_443;
	wire [0 : 0] fresh_wire_444;
	wire [0 : 0] fresh_wire_445;
	wire [0 : 0] fresh_wire_446;
	wire [0 : 0] fresh_wire_447;
	wire [0 : 0] fresh_wire_448;
	wire [0 : 0] fresh_wire_449;
	wire [0 : 0] fresh_wire_450;
	wire [0 : 0] fresh_wire_451;
	wire [0 : 0] fresh_wire_452;
	wire [0 : 0] fresh_wire_453;
	wire [0 : 0] fresh_wire_454;
	wire [0 : 0] fresh_wire_455;
	wire [0 : 0] fresh_wire_456;
	wire [15 : 0] fresh_wire_457;
	wire [15 : 0] fresh_wire_458;
	wire [15 : 0] fresh_wire_459;
	wire [0 : 0] fresh_wire_460;
	wire [15 : 0] fresh_wire_461;
	wire [15 : 0] fresh_wire_462;
	wire [15 : 0] fresh_wire_463;
	wire [0 : 0] fresh_wire_464;
	wire [15 : 0] fresh_wire_465;
	wire [15 : 0] fresh_wire_466;
	wire [15 : 0] fresh_wire_467;
	wire [0 : 0] fresh_wire_468;
	wire [15 : 0] fresh_wire_469;
	wire [15 : 0] fresh_wire_470;
	wire [15 : 0] fresh_wire_471;
	wire [0 : 0] fresh_wire_472;
	wire [1 : 0] fresh_wire_473;
	wire [1 : 0] fresh_wire_474;
	wire [1 : 0] fresh_wire_475;
	wire [0 : 0] fresh_wire_476;
	wire [1 : 0] fresh_wire_477;
	wire [1 : 0] fresh_wire_478;
	wire [1 : 0] fresh_wire_479;
	wire [0 : 0] fresh_wire_480;
	wire [1 : 0] fresh_wire_481;
	wire [1 : 0] fresh_wire_482;
	wire [1 : 0] fresh_wire_483;
	wire [0 : 0] fresh_wire_484;
	wire [1 : 0] fresh_wire_485;
	wire [1 : 0] fresh_wire_486;
	wire [1 : 0] fresh_wire_487;
	wire [0 : 0] fresh_wire_488;
	wire [1 : 0] fresh_wire_489;
	wire [1 : 0] fresh_wire_490;
	wire [1 : 0] fresh_wire_491;
	wire [0 : 0] fresh_wire_492;
	wire [1 : 0] fresh_wire_493;
	wire [1 : 0] fresh_wire_494;
	wire [1 : 0] fresh_wire_495;
	wire [0 : 0] fresh_wire_496;
	wire [0 : 0] fresh_wire_497;
	wire [0 : 0] fresh_wire_498;
	wire [0 : 0] fresh_wire_499;
	wire [0 : 0] fresh_wire_500;
	wire [0 : 0] fresh_wire_501;
	wire [0 : 0] fresh_wire_502;
	wire [0 : 0] fresh_wire_503;
	wire [0 : 0] fresh_wire_504;
	wire [0 : 0] fresh_wire_505;
	wire [0 : 0] fresh_wire_506;
	wire [0 : 0] fresh_wire_507;
	wire [0 : 0] fresh_wire_508;
	wire [0 : 0] fresh_wire_509;
	wire [0 : 0] fresh_wire_510;
	wire [0 : 0] fresh_wire_511;
	wire [0 : 0] fresh_wire_512;
	wire [0 : 0] fresh_wire_513;
	wire [0 : 0] fresh_wire_514;
	wire [0 : 0] fresh_wire_515;
	wire [0 : 0] fresh_wire_516;
	wire [0 : 0] fresh_wire_517;
	wire [0 : 0] fresh_wire_518;
	wire [0 : 0] fresh_wire_519;
	wire [0 : 0] fresh_wire_520;
	wire [0 : 0] fresh_wire_521;
	wire [0 : 0] fresh_wire_522;
	wire [0 : 0] fresh_wire_523;
	wire [0 : 0] fresh_wire_524;
	wire [0 : 0] fresh_wire_525;
	wire [0 : 0] fresh_wire_526;
	wire [0 : 0] fresh_wire_527;
	wire [0 : 0] fresh_wire_528;
	wire [0 : 0] fresh_wire_529;
	wire [0 : 0] fresh_wire_530;
	wire [0 : 0] fresh_wire_531;
	wire [0 : 0] fresh_wire_532;
	wire [0 : 0] fresh_wire_533;
	wire [0 : 0] fresh_wire_534;
	wire [0 : 0] fresh_wire_535;
	wire [0 : 0] fresh_wire_536;
	wire [15 : 0] fresh_wire_537;
	wire [15 : 0] fresh_wire_538;
	wire [15 : 0] fresh_wire_539;
	wire [0 : 0] fresh_wire_540;
	wire [15 : 0] fresh_wire_541;
	wire [15 : 0] fresh_wire_542;
	wire [15 : 0] fresh_wire_543;
	wire [0 : 0] fresh_wire_544;
	wire [15 : 0] fresh_wire_545;
	wire [15 : 0] fresh_wire_546;
	wire [15 : 0] fresh_wire_547;
	wire [0 : 0] fresh_wire_548;
	wire [15 : 0] fresh_wire_549;
	wire [15 : 0] fresh_wire_550;
	wire [15 : 0] fresh_wire_551;
	wire [0 : 0] fresh_wire_552;
	wire [15 : 0] fresh_wire_553;
	wire [15 : 0] fresh_wire_554;
	wire [15 : 0] fresh_wire_555;
	wire [0 : 0] fresh_wire_556;
	wire [15 : 0] fresh_wire_557;
	wire [15 : 0] fresh_wire_558;
	wire [15 : 0] fresh_wire_559;
	wire [0 : 0] fresh_wire_560;
	wire [15 : 0] fresh_wire_561;
	wire [15 : 0] fresh_wire_562;
	wire [15 : 0] fresh_wire_563;
	wire [0 : 0] fresh_wire_564;
	wire [15 : 0] fresh_wire_565;
	wire [15 : 0] fresh_wire_566;
	wire [15 : 0] fresh_wire_567;
	wire [0 : 0] fresh_wire_568;
	wire [15 : 0] fresh_wire_569;
	wire [15 : 0] fresh_wire_570;
	wire [15 : 0] fresh_wire_571;
	wire [0 : 0] fresh_wire_572;
	wire [0 : 0] fresh_wire_573;
	wire [0 : 0] fresh_wire_574;
	wire [0 : 0] fresh_wire_575;
	wire [0 : 0] fresh_wire_576;
	wire [0 : 0] fresh_wire_577;
	wire [0 : 0] fresh_wire_578;
	wire [0 : 0] fresh_wire_579;
	wire [0 : 0] fresh_wire_580;
	wire [0 : 0] fresh_wire_581;
	wire [0 : 0] fresh_wire_582;
	wire [0 : 0] fresh_wire_583;
	wire [0 : 0] fresh_wire_584;
	wire [0 : 0] fresh_wire_585;
	wire [0 : 0] fresh_wire_586;
	wire [0 : 0] fresh_wire_587;
	wire [0 : 0] fresh_wire_588;
	wire [0 : 0] fresh_wire_589;
	wire [0 : 0] fresh_wire_590;
	wire [0 : 0] fresh_wire_591;
	wire [0 : 0] fresh_wire_592;
	wire [15 : 0] fresh_wire_593;
	wire [31 : 0] fresh_wire_594;
	wire [31 : 0] fresh_wire_595;
	wire [31 : 0] fresh_wire_596;
	wire [31 : 0] fresh_wire_597;
	wire [31 : 0] fresh_wire_598;
	wire [31 : 0] fresh_wire_599;
	wire [31 : 0] fresh_wire_600;
	wire [0 : 0] fresh_wire_601;
	wire [15 : 0] fresh_wire_602;
	wire [15 : 0] fresh_wire_603;
	wire [15 : 0] fresh_wire_604;
	wire [0 : 0] fresh_wire_605;
	wire [0 : 0] fresh_wire_606;
	wire [15 : 0] fresh_wire_607;
	wire [15 : 0] fresh_wire_608;
	wire [15 : 0] fresh_wire_609;
	wire [0 : 0] fresh_wire_610;
	wire [1 : 0] fresh_wire_611;
	wire [1 : 0] fresh_wire_612;
	wire [1 : 0] fresh_wire_613;
	wire [0 : 0] fresh_wire_614;
	wire [0 : 0] fresh_wire_615;
	wire [0 : 0] fresh_wire_616;
	wire [0 : 0] fresh_wire_617;
	wire [0 : 0] fresh_wire_618;
	wire [0 : 0] fresh_wire_619;
	wire [0 : 0] fresh_wire_620;
	wire [0 : 0] fresh_wire_621;
	wire [0 : 0] fresh_wire_622;
	wire [1 : 0] fresh_wire_623;
	wire [1 : 0] fresh_wire_624;
	wire [0 : 0] fresh_wire_625;
	wire [1 : 0] fresh_wire_626;
	wire [1 : 0] fresh_wire_627;
	wire [0 : 0] fresh_wire_628;
	wire [0 : 0] fresh_wire_629;
	wire [0 : 0] fresh_wire_630;
	wire [0 : 0] fresh_wire_631;
	wire [1 : 0] fresh_wire_632;
	wire [1 : 0] fresh_wire_633;
	wire [0 : 0] fresh_wire_634;
	wire [1 : 0] fresh_wire_635;
	wire [1 : 0] fresh_wire_636;
	wire [0 : 0] fresh_wire_637;
	wire [0 : 0] fresh_wire_638;
	wire [0 : 0] fresh_wire_639;
	wire [0 : 0] fresh_wire_640;
	wire [0 : 0] fresh_wire_641;
	wire [0 : 0] fresh_wire_642;
	wire [0 : 0] fresh_wire_643;
	wire [0 : 0] fresh_wire_644;
	wire [0 : 0] fresh_wire_645;
	wire [0 : 0] fresh_wire_646;
	wire [0 : 0] fresh_wire_647;
	wire [0 : 0] fresh_wire_648;
	wire [0 : 0] fresh_wire_649;
	wire [0 : 0] fresh_wire_650;
	wire [0 : 0] fresh_wire_651;
	wire [0 : 0] fresh_wire_652;
	wire [0 : 0] fresh_wire_653;
	wire [0 : 0] fresh_wire_654;
	wire [0 : 0] fresh_wire_655;
	wire [0 : 0] fresh_wire_656;
	wire [0 : 0] fresh_wire_657;
	wire [0 : 0] fresh_wire_658;
	wire [0 : 0] fresh_wire_659;
	wire [0 : 0] fresh_wire_660;
	wire [0 : 0] fresh_wire_661;
	wire [0 : 0] fresh_wire_662;
	wire [0 : 0] fresh_wire_663;
	wire [0 : 0] fresh_wire_664;
	wire [1 : 0] fresh_wire_665;
	wire [1 : 0] fresh_wire_666;
	wire [0 : 0] fresh_wire_667;
	wire [0 : 0] fresh_wire_668;
	wire [47 : 0] fresh_wire_669;
	wire [47 : 0] fresh_wire_670;
	wire [0 : 0] fresh_wire_671;
	wire [0 : 0] fresh_wire_672;
	wire [0 : 0] fresh_wire_673;
	wire [0 : 0] fresh_wire_674;
	wire [0 : 0] fresh_wire_675;
	wire [0 : 0] fresh_wire_676;
	wire [0 : 0] fresh_wire_677;
	wire [0 : 0] fresh_wire_678;
	wire [0 : 0] fresh_wire_679;
	wire [1 : 0] fresh_wire_680;
	wire [1 : 0] fresh_wire_681;
	wire [1 : 0] fresh_wire_682;
	wire [0 : 0] fresh_wire_683;
	wire [1 : 0] fresh_wire_684;
	wire [1 : 0] fresh_wire_685;
	wire [1 : 0] fresh_wire_686;
	wire [0 : 0] fresh_wire_687;
	wire [31 : 0] fresh_wire_688;
	wire [31 : 0] fresh_wire_689;
	wire [31 : 0] fresh_wire_690;
	wire [0 : 0] fresh_wire_691;
	wire [31 : 0] fresh_wire_692;
	wire [31 : 0] fresh_wire_693;
	wire [31 : 0] fresh_wire_694;
	wire [0 : 0] fresh_wire_695;
	wire [31 : 0] fresh_wire_696;
	wire [31 : 0] fresh_wire_697;
	wire [31 : 0] fresh_wire_698;
	wire [0 : 0] fresh_wire_699;
	wire [31 : 0] fresh_wire_700;
	wire [31 : 0] fresh_wire_701;
	wire [31 : 0] fresh_wire_702;
	wire [0 : 0] fresh_wire_703;
	wire [31 : 0] fresh_wire_704;
	wire [31 : 0] fresh_wire_705;
	wire [31 : 0] fresh_wire_706;
	wire [0 : 0] fresh_wire_707;
	wire [31 : 0] fresh_wire_708;
	wire [31 : 0] fresh_wire_709;
	wire [31 : 0] fresh_wire_710;
	wire [0 : 0] fresh_wire_711;
	wire [31 : 0] fresh_wire_712;
	wire [31 : 0] fresh_wire_713;
	wire [31 : 0] fresh_wire_714;
	wire [0 : 0] fresh_wire_715;
	wire [1 : 0] fresh_wire_716;
	wire [1 : 0] fresh_wire_717;
	wire [1 : 0] fresh_wire_718;
	wire [0 : 0] fresh_wire_719;
	wire [1 : 0] fresh_wire_720;
	wire [1 : 0] fresh_wire_721;
	wire [1 : 0] fresh_wire_722;
	wire [1 : 0] fresh_wire_723;
	wire [1 : 0] fresh_wire_724;
	wire [1 : 0] fresh_wire_725;
	wire [0 : 0] fresh_wire_726;
	wire [0 : 0] fresh_wire_727;
	wire [0 : 0] fresh_wire_728;
	wire [0 : 0] fresh_wire_729;
	wire [0 : 0] fresh_wire_730;
	wire [0 : 0] fresh_wire_731;
	wire [0 : 0] fresh_wire_732;
	wire [0 : 0] fresh_wire_733;
	wire [0 : 0] fresh_wire_734;
	wire [0 : 0] fresh_wire_735;
	wire [0 : 0] fresh_wire_736;
	wire [0 : 0] fresh_wire_737;
	wire [0 : 0] fresh_wire_738;
	wire [0 : 0] fresh_wire_739;
	wire [0 : 0] fresh_wire_740;
	wire [0 : 0] fresh_wire_741;
	wire [0 : 0] fresh_wire_742;
	wire [0 : 0] fresh_wire_743;
	wire [1 : 0] fresh_wire_744;
	wire [1 : 0] fresh_wire_745;
	wire [0 : 0] fresh_wire_746;
	wire [1 : 0] fresh_wire_747;
	wire [1 : 0] fresh_wire_748;
	wire [0 : 0] fresh_wire_749;
	wire [1 : 0] fresh_wire_750;
	wire [1 : 0] fresh_wire_751;
	wire [0 : 0] fresh_wire_752;
	wire [1 : 0] fresh_wire_753;
	wire [1 : 0] fresh_wire_754;
	wire [0 : 0] fresh_wire_755;
	wire [1 : 0] fresh_wire_756;
	wire [1 : 0] fresh_wire_757;
	wire [0 : 0] fresh_wire_758;
	wire [0 : 0] fresh_wire_759;
	wire [0 : 0] fresh_wire_760;
	wire [0 : 0] fresh_wire_761;
	wire [0 : 0] fresh_wire_762;
	wire [0 : 0] fresh_wire_763;
	wire [0 : 0] fresh_wire_764;
	wire [0 : 0] fresh_wire_765;
	wire [0 : 0] fresh_wire_766;
	wire [0 : 0] fresh_wire_767;
	wire [0 : 0] fresh_wire_768;
	wire [0 : 0] fresh_wire_769;
	wire [0 : 0] fresh_wire_770;
	wire [0 : 0] fresh_wire_771;
	wire [0 : 0] fresh_wire_772;
	wire [0 : 0] fresh_wire_773;
	wire [0 : 0] fresh_wire_774;
	wire [0 : 0] fresh_wire_775;
	wire [0 : 0] fresh_wire_776;
	wire [0 : 0] fresh_wire_777;
	wire [0 : 0] fresh_wire_778;
	wire [0 : 0] fresh_wire_779;
	wire [0 : 0] fresh_wire_780;
	wire [0 : 0] fresh_wire_781;
	wire [0 : 0] fresh_wire_782;
	wire [0 : 0] fresh_wire_783;
	wire [0 : 0] fresh_wire_784;
	wire [0 : 0] fresh_wire_785;
	wire [0 : 0] fresh_wire_786;
	wire [0 : 0] fresh_wire_787;
	wire [0 : 0] fresh_wire_788;
	wire [0 : 0] fresh_wire_789;
	wire [0 : 0] fresh_wire_790;
	wire [0 : 0] fresh_wire_791;
	wire [0 : 0] fresh_wire_792;
	wire [0 : 0] fresh_wire_793;
	wire [0 : 0] fresh_wire_794;
	wire [0 : 0] fresh_wire_795;
	wire [0 : 0] fresh_wire_796;
	wire [0 : 0] fresh_wire_797;
	wire [0 : 0] fresh_wire_798;
	wire [0 : 0] fresh_wire_799;
	wire [0 : 0] fresh_wire_800;
	wire [0 : 0] fresh_wire_801;
	wire [0 : 0] fresh_wire_802;
	wire [0 : 0] fresh_wire_803;
	wire [0 : 0] fresh_wire_804;
	wire [0 : 0] fresh_wire_805;
	wire [0 : 0] fresh_wire_806;
	wire [0 : 0] fresh_wire_807;
	wire [0 : 0] fresh_wire_808;
	wire [0 : 0] fresh_wire_809;
	wire [0 : 0] fresh_wire_810;
	wire [0 : 0] fresh_wire_811;
	wire [0 : 0] fresh_wire_812;
	wire [0 : 0] fresh_wire_813;
	wire [0 : 0] fresh_wire_814;
	wire [0 : 0] fresh_wire_815;
	wire [0 : 0] fresh_wire_816;
	wire [0 : 0] fresh_wire_817;
	wire [0 : 0] fresh_wire_818;
	wire [0 : 0] fresh_wire_819;
	wire [0 : 0] fresh_wire_820;
	wire [0 : 0] fresh_wire_821;
	wire [0 : 0] fresh_wire_822;
	wire [0 : 0] fresh_wire_823;
	wire [0 : 0] fresh_wire_824;
	wire [0 : 0] fresh_wire_825;
	wire [0 : 0] fresh_wire_826;
	wire [0 : 0] fresh_wire_827;
	wire [0 : 0] fresh_wire_828;
	wire [0 : 0] fresh_wire_829;
	wire [0 : 0] fresh_wire_830;
	wire [0 : 0] fresh_wire_831;
	wire [0 : 0] fresh_wire_832;
	wire [0 : 0] fresh_wire_833;
	wire [0 : 0] fresh_wire_834;
	wire [0 : 0] fresh_wire_835;
	wire [0 : 0] fresh_wire_836;
	wire [0 : 0] fresh_wire_837;
	wire [0 : 0] fresh_wire_838;
	wire [0 : 0] fresh_wire_839;
	wire [0 : 0] fresh_wire_840;
	wire [0 : 0] fresh_wire_841;
	wire [0 : 0] fresh_wire_842;
	wire [0 : 0] fresh_wire_843;
	wire [0 : 0] fresh_wire_844;
	wire [0 : 0] fresh_wire_845;
	wire [0 : 0] fresh_wire_846;
	wire [0 : 0] fresh_wire_847;
	wire [0 : 0] fresh_wire_848;
	wire [0 : 0] fresh_wire_849;
	wire [0 : 0] fresh_wire_850;
	wire [0 : 0] fresh_wire_851;
	wire [0 : 0] fresh_wire_852;
	wire [0 : 0] fresh_wire_853;
	wire [0 : 0] fresh_wire_854;
	wire [0 : 0] fresh_wire_855;
	wire [0 : 0] fresh_wire_856;
	wire [1 : 0] fresh_wire_857;
	wire [1 : 0] fresh_wire_858;
	wire [0 : 0] fresh_wire_859;
	wire [0 : 0] fresh_wire_860;
	wire [47 : 0] fresh_wire_861;
	wire [47 : 0] fresh_wire_862;
	wire [0 : 0] fresh_wire_863;
	wire [15 : 0] fresh_wire_864;
	wire [15 : 0] fresh_wire_865;
	wire [15 : 0] fresh_wire_866;
	wire [0 : 0] fresh_wire_867;
	wire [15 : 0] fresh_wire_868;
	wire [15 : 0] fresh_wire_869;
	wire [15 : 0] fresh_wire_870;
	wire [0 : 0] fresh_wire_871;
	wire [15 : 0] fresh_wire_872;
	wire [15 : 0] fresh_wire_873;
	wire [15 : 0] fresh_wire_874;
	wire [0 : 0] fresh_wire_875;
	wire [15 : 0] fresh_wire_876;
	wire [15 : 0] fresh_wire_877;
	wire [15 : 0] fresh_wire_878;
	wire [0 : 0] fresh_wire_879;
	wire [0 : 0] fresh_wire_880;
	wire [0 : 0] fresh_wire_881;
	wire [0 : 0] fresh_wire_882;
	wire [0 : 0] fresh_wire_883;
	wire [0 : 0] fresh_wire_884;
	wire [0 : 0] fresh_wire_885;
	wire [0 : 0] fresh_wire_886;
	wire [0 : 0] fresh_wire_887;
	wire [0 : 0] fresh_wire_888;
	wire [0 : 0] fresh_wire_889;
	wire [0 : 0] fresh_wire_890;
	wire [0 : 0] fresh_wire_891;
	wire [0 : 0] fresh_wire_892;
	wire [0 : 0] fresh_wire_893;
	wire [0 : 0] fresh_wire_894;
	wire [0 : 0] fresh_wire_895;
	wire [1 : 0] fresh_wire_896;
	wire [1 : 0] fresh_wire_897;
	wire [1 : 0] fresh_wire_898;
	wire [0 : 0] fresh_wire_899;
	wire [1 : 0] fresh_wire_900;
	wire [1 : 0] fresh_wire_901;
	wire [1 : 0] fresh_wire_902;
	wire [0 : 0] fresh_wire_903;
	wire [1 : 0] fresh_wire_904;
	wire [1 : 0] fresh_wire_905;
	wire [1 : 0] fresh_wire_906;
	wire [0 : 0] fresh_wire_907;
	wire [1 : 0] fresh_wire_908;
	wire [1 : 0] fresh_wire_909;
	wire [1 : 0] fresh_wire_910;
	wire [0 : 0] fresh_wire_911;
	wire [1 : 0] fresh_wire_912;
	wire [1 : 0] fresh_wire_913;
	wire [1 : 0] fresh_wire_914;
	wire [0 : 0] fresh_wire_915;
	wire [47 : 0] fresh_wire_916;
	wire [47 : 0] fresh_wire_917;
	wire [47 : 0] fresh_wire_918;
	wire [0 : 0] fresh_wire_919;
	wire [47 : 0] fresh_wire_920;
	wire [47 : 0] fresh_wire_921;
	wire [47 : 0] fresh_wire_922;
	wire [0 : 0] fresh_wire_923;
	wire [1 : 0] fresh_wire_924;
	wire [1 : 0] fresh_wire_925;
	wire [1 : 0] fresh_wire_926;
	wire [0 : 0] fresh_wire_927;
	wire [0 : 0] fresh_wire_928;
	wire [0 : 0] fresh_wire_929;
	wire [0 : 0] fresh_wire_930;
	wire [0 : 0] fresh_wire_931;
	wire [0 : 0] fresh_wire_932;
	wire [0 : 0] fresh_wire_933;
	wire [0 : 0] fresh_wire_934;
	wire [0 : 0] fresh_wire_935;
	wire [0 : 0] fresh_wire_936;
	wire [0 : 0] fresh_wire_937;
	wire [15 : 0] fresh_wire_938;
	wire [15 : 0] fresh_wire_939;
	wire [0 : 0] fresh_wire_940;
	wire [15 : 0] fresh_wire_941;
	wire [15 : 0] fresh_wire_942;
	wire [15 : 0] fresh_wire_943;
	wire [0 : 0] fresh_wire_944;
	wire [15 : 0] fresh_wire_945;
	wire [15 : 0] fresh_wire_946;
	wire [15 : 0] fresh_wire_947;
	wire [0 : 0] fresh_wire_948;
	wire [0 : 0] fresh_wire_949;
	wire [15 : 0] fresh_wire_950;
	wire [15 : 0] fresh_wire_951;
	wire [15 : 0] fresh_wire_952;
	wire [0 : 0] fresh_wire_953;
	wire [15 : 0] fresh_wire_954;
	wire [15 : 0] fresh_wire_955;
	wire [15 : 0] fresh_wire_956;
	wire [0 : 0] fresh_wire_957;
	wire [0 : 0] fresh_wire_958;
	wire [0 : 0] fresh_wire_959;
	wire [0 : 0] fresh_wire_960;
	wire [0 : 0] fresh_wire_961;
	wire [0 : 0] fresh_wire_962;
	wire [0 : 0] fresh_wire_963;
	wire [0 : 0] fresh_wire_964;
	wire [0 : 0] fresh_wire_965;
	wire [0 : 0] fresh_wire_966;
	wire [0 : 0] fresh_wire_967;
	wire [0 : 0] fresh_wire_968;
	wire [0 : 0] fresh_wire_969;
	wire [0 : 0] fresh_wire_970;
	wire [0 : 0] fresh_wire_971;
	wire [0 : 0] fresh_wire_972;
	wire [0 : 0] fresh_wire_973;
	wire [15 : 0] fresh_wire_974;
	wire [15 : 0] fresh_wire_975;
	wire [15 : 0] fresh_wire_976;
	wire [0 : 0] fresh_wire_977;
	wire [0 : 0] fresh_wire_978;
	wire [0 : 0] fresh_wire_979;
	wire [0 : 0] fresh_wire_980;
	wire [0 : 0] fresh_wire_981;
	wire [0 : 0] fresh_wire_982;
	wire [0 : 0] fresh_wire_983;
	wire [0 : 0] fresh_wire_984;
	wire [0 : 0] fresh_wire_985;
	wire [0 : 0] fresh_wire_986;
	wire [0 : 0] fresh_wire_987;
	wire [0 : 0] fresh_wire_988;
	wire [0 : 0] fresh_wire_989;
	wire [0 : 0] fresh_wire_990;
	wire [0 : 0] fresh_wire_991;
	wire [0 : 0] fresh_wire_992;
	wire [0 : 0] fresh_wire_993;
	wire [8 : 0] fresh_wire_994;
	wire [8 : 0] fresh_wire_995;
	wire [8 : 0] fresh_wire_996;
	wire [0 : 0] fresh_wire_997;
	wire [0 : 0] fresh_wire_998;
	wire [0 : 0] fresh_wire_999;
	wire [0 : 0] fresh_wire_1000;
	wire [0 : 0] fresh_wire_1001;
	wire [0 : 0] fresh_wire_1002;
	wire [0 : 0] fresh_wire_1003;
	wire [0 : 0] fresh_wire_1004;
	wire [0 : 0] fresh_wire_1005;
	wire [0 : 0] fresh_wire_1006;
	wire [8 : 0] fresh_wire_1007;
	wire [8 : 0] fresh_wire_1008;
	wire [8 : 0] fresh_wire_1009;
	wire [0 : 0] fresh_wire_1010;
	wire [0 : 0] fresh_wire_1011;
	wire [0 : 0] fresh_wire_1012;
	wire [0 : 0] fresh_wire_1013;
	wire [0 : 0] fresh_wire_1014;
	wire [0 : 0] fresh_wire_1015;
	wire [0 : 0] fresh_wire_1016;
	wire [0 : 0] fresh_wire_1017;
	wire [0 : 0] fresh_wire_1018;
	wire [0 : 0] fresh_wire_1019;
	wire [0 : 0] fresh_wire_1020;
	wire [8 : 0] fresh_wire_1021;
	wire [15 : 0] fresh_wire_1022;
	wire [8 : 0] fresh_wire_1023;
	wire [15 : 0] fresh_wire_1024;
	wire [0 : 0] fresh_wire_1025;
	wire [0 : 0] fresh_wire_1026;
	wire [0 : 0] fresh_wire_1027;
	wire [0 : 0] fresh_wire_1028;
	wire [0 : 0] fresh_wire_1029;
	wire [0 : 0] fresh_wire_1030;
	wire [0 : 0] fresh_wire_1031;
	wire [0 : 0] fresh_wire_1032;
	wire [0 : 0] fresh_wire_1033;
	wire [0 : 0] fresh_wire_1034;
	wire [0 : 0] fresh_wire_1035;
	wire [15 : 0] fresh_wire_1036;
	wire [15 : 0] fresh_wire_1037;
	wire [0 : 0] fresh_wire_1038;
	wire [15 : 0] fresh_wire_1039;
	wire [15 : 0] fresh_wire_1040;
	wire [15 : 0] fresh_wire_1041;
	wire [0 : 0] fresh_wire_1042;
	wire [15 : 0] fresh_wire_1043;
	wire [15 : 0] fresh_wire_1044;
	wire [15 : 0] fresh_wire_1045;
	wire [0 : 0] fresh_wire_1046;
	wire [0 : 0] fresh_wire_1047;
	wire [15 : 0] fresh_wire_1048;
	wire [15 : 0] fresh_wire_1049;
	wire [15 : 0] fresh_wire_1050;
	wire [0 : 0] fresh_wire_1051;
	wire [15 : 0] fresh_wire_1052;
	wire [15 : 0] fresh_wire_1053;
	wire [15 : 0] fresh_wire_1054;
	wire [0 : 0] fresh_wire_1055;
	wire [0 : 0] fresh_wire_1056;
	wire [0 : 0] fresh_wire_1057;
	wire [0 : 0] fresh_wire_1058;
	wire [0 : 0] fresh_wire_1059;
	wire [0 : 0] fresh_wire_1060;
	wire [0 : 0] fresh_wire_1061;
	wire [0 : 0] fresh_wire_1062;
	wire [0 : 0] fresh_wire_1063;
	wire [0 : 0] fresh_wire_1064;
	wire [0 : 0] fresh_wire_1065;
	wire [0 : 0] fresh_wire_1066;
	wire [0 : 0] fresh_wire_1067;
	wire [0 : 0] fresh_wire_1068;
	wire [0 : 0] fresh_wire_1069;
	wire [0 : 0] fresh_wire_1070;
	wire [0 : 0] fresh_wire_1071;
	wire [15 : 0] fresh_wire_1072;
	wire [15 : 0] fresh_wire_1073;
	wire [15 : 0] fresh_wire_1074;
	wire [0 : 0] fresh_wire_1075;
	wire [0 : 0] fresh_wire_1076;
	wire [0 : 0] fresh_wire_1077;
	wire [0 : 0] fresh_wire_1078;
	wire [0 : 0] fresh_wire_1079;
	wire [0 : 0] fresh_wire_1080;
	wire [0 : 0] fresh_wire_1081;
	wire [0 : 0] fresh_wire_1082;
	wire [0 : 0] fresh_wire_1083;
	wire [0 : 0] fresh_wire_1084;
	wire [0 : 0] fresh_wire_1085;
	wire [0 : 0] fresh_wire_1086;
	wire [0 : 0] fresh_wire_1087;
	wire [0 : 0] fresh_wire_1088;
	wire [0 : 0] fresh_wire_1089;
	wire [0 : 0] fresh_wire_1090;
	wire [0 : 0] fresh_wire_1091;
	wire [8 : 0] fresh_wire_1092;
	wire [8 : 0] fresh_wire_1093;
	wire [8 : 0] fresh_wire_1094;
	wire [0 : 0] fresh_wire_1095;
	wire [0 : 0] fresh_wire_1096;
	wire [0 : 0] fresh_wire_1097;
	wire [0 : 0] fresh_wire_1098;
	wire [0 : 0] fresh_wire_1099;
	wire [0 : 0] fresh_wire_1100;
	wire [0 : 0] fresh_wire_1101;
	wire [0 : 0] fresh_wire_1102;
	wire [0 : 0] fresh_wire_1103;
	wire [0 : 0] fresh_wire_1104;
	wire [8 : 0] fresh_wire_1105;
	wire [8 : 0] fresh_wire_1106;
	wire [8 : 0] fresh_wire_1107;
	wire [0 : 0] fresh_wire_1108;
	wire [0 : 0] fresh_wire_1109;
	wire [0 : 0] fresh_wire_1110;
	wire [0 : 0] fresh_wire_1111;
	wire [0 : 0] fresh_wire_1112;
	wire [0 : 0] fresh_wire_1113;
	wire [0 : 0] fresh_wire_1114;
	wire [0 : 0] fresh_wire_1115;
	wire [0 : 0] fresh_wire_1116;
	wire [0 : 0] fresh_wire_1117;
	wire [0 : 0] fresh_wire_1118;
	wire [8 : 0] fresh_wire_1119;
	wire [15 : 0] fresh_wire_1120;
	wire [8 : 0] fresh_wire_1121;
	wire [15 : 0] fresh_wire_1122;
	wire [0 : 0] fresh_wire_1123;
	wire [16 : 0] fresh_wire_1124;
	wire [33 : 0] fresh_wire_1125;
	wire [33 : 0] fresh_wire_1126;
	wire [33 : 0] fresh_wire_1127;
	wire [33 : 0] fresh_wire_1128;
	wire [15 : 0] fresh_wire_1129;
	wire [16 : 0] fresh_wire_1130;
	wire [16 : 0] fresh_wire_1131;
	wire [16 : 0] fresh_wire_1132;
	wire [16 : 0] fresh_wire_1133;
	wire [16 : 0] fresh_wire_1134;
	wire [16 : 0] fresh_wire_1135;
	wire [16 : 0] fresh_wire_1136;
	wire [16 : 0] fresh_wire_1137;
	wire [33 : 0] fresh_wire_1138;
	wire [33 : 0] fresh_wire_1139;
	wire [33 : 0] fresh_wire_1140;
	wire [33 : 0] fresh_wire_1141;
	wire [15 : 0] fresh_wire_1142;
	wire [16 : 0] fresh_wire_1143;
	wire [15 : 0] fresh_wire_1144;
	wire [16 : 0] fresh_wire_1145;
	wire [16 : 0] fresh_wire_1146;
	wire [16 : 0] fresh_wire_1147;
	wire [16 : 0] fresh_wire_1148;
	wire [16 : 0] fresh_wire_1149;
	wire [16 : 0] fresh_wire_1150;
	wire [16 : 0] fresh_wire_1151;
	wire [0 : 0] fresh_wire_1152;
	wire [0 : 0] fresh_wire_1153;
	wire [15 : 0] fresh_wire_1154;
	wire [15 : 0] fresh_wire_1155;
	wire [15 : 0] fresh_wire_1156;
	wire [15 : 0] fresh_wire_1157;
	wire [15 : 0] fresh_wire_1158;
	wire [15 : 0] fresh_wire_1159;
	wire [15 : 0] fresh_wire_1160;
	wire [15 : 0] fresh_wire_1161;
	wire [15 : 0] fresh_wire_1162;
	wire [0 : 0] fresh_wire_1163;
	wire [33 : 0] fresh_wire_1164;
	wire [16 : 0] fresh_wire_1165;
	wire [16 : 0] fresh_wire_1166;
	wire [0 : 0] fresh_wire_1167;
	wire [33 : 0] fresh_wire_1168;
	wire [0 : 0] fresh_wire_1169;
	wire [0 : 0] fresh_wire_1170;
	wire [0 : 0] fresh_wire_1171;
	wire [0 : 0] fresh_wire_1172;
	wire [0 : 0] fresh_wire_1173;
	wire [16 : 0] fresh_wire_1174;
	wire [0 : 0] fresh_wire_1175;
	wire [0 : 0] fresh_wire_1176;
	wire [0 : 0] fresh_wire_1177;
	wire [0 : 0] fresh_wire_1178;
	wire [0 : 0] fresh_wire_1179;
	wire [0 : 0] fresh_wire_1180;
	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) aux_div_pad_port_cell(.PORT_ID_IN(fresh_wire_0),
.PORT_ID_OUT(aux_div_pad));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) cell_149_const_replacement(.PORT_ID_OUT(fresh_wire_1153));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) cell_261940_const_replacement(.PORT_ID_OUT(fresh_wire_1163));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(34'h000000007),
.PARAM_WIDTH(32'h00000022)) cell_261945_const_replacement(.PORT_ID_OUT(fresh_wire_1164));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(16'h0001),
.PARAM_WIDTH(32'h00000010)) cell_26382_const_replacement(.PORT_ID_OUT(fresh_wire_1154));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(16'h0002),
.PARAM_WIDTH(32'h00000010)) cell_26400_const_replacement(.PORT_ID_OUT(fresh_wire_1155));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(16'h0002),
.PARAM_WIDTH(32'h00000010)) cell_26409_const_replacement(.PORT_ID_OUT(fresh_wire_1156));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(16'h0001),
.PARAM_WIDTH(32'h00000010)) cell_26415_const_replacement(.PORT_ID_OUT(fresh_wire_1157));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(17'h00000),
.PARAM_WIDTH(32'h00000011)) cell_264252_const_replacement(.PORT_ID_OUT(fresh_wire_1166));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(17'h00000),
.PARAM_WIDTH(32'h00000011)) cell_264255_const_replacement(.PORT_ID_OUT(fresh_wire_1165));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(16'h000a),
.PARAM_WIDTH(32'h00000010)) cell_26436_const_replacement(.PORT_ID_OUT(fresh_wire_1158));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(16'h000a),
.PARAM_WIDTH(32'h00000010)) cell_26550_const_replacement(.PORT_ID_OUT(fresh_wire_1159));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_26608_const_replacement(.PORT_ID_OUT(fresh_wire_1175));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_26618_const_replacement(.PORT_ID_OUT(fresh_wire_1176));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_26641_const_replacement(.PORT_ID_OUT(fresh_wire_1177));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_26648_const_replacement(.PORT_ID_OUT(fresh_wire_1178));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_26668_const_replacement(.PORT_ID_OUT(fresh_wire_1179));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) cell_26671_const_replacement(.PORT_ID_OUT(fresh_wire_1180));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) cell_267321_const_replacement(.PORT_ID_OUT(fresh_wire_1167));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(34'h000000007),
.PARAM_WIDTH(32'h00000022)) cell_267326_const_replacement(.PORT_ID_OUT(fresh_wire_1168));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(16'h000a),
.PARAM_WIDTH(32'h00000010)) cell_26849_const_replacement(.PORT_ID_OUT(fresh_wire_1160));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(16'h0004),
.PARAM_WIDTH(32'h00000010)) cell_26860_const_replacement(.PORT_ID_OUT(fresh_wire_1161));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(16'h0005),
.PARAM_WIDTH(32'h00000010)) cell_26866_const_replacement(.PORT_ID_OUT(fresh_wire_1162));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_269371_const_replacement(.PORT_ID_OUT(fresh_wire_1169));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_27034_const_replacement(.PORT_ID_OUT(fresh_wire_1170));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_27039_const_replacement(.PORT_ID_OUT(fresh_wire_1171));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_27064_const_replacement(.PORT_ID_OUT(fresh_wire_1172));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_27069_const_replacement(.PORT_ID_OUT(fresh_wire_1173));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(17'h00000),
.PARAM_WIDTH(32'h00000011)) cell_296571_const_replacement(.PORT_ID_OUT(fresh_wire_1174));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) clk_ext_in_port_cell(.PORT_ID_IN(clk_ext_in),
.PORT_ID_OUT(fresh_wire_1));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) clk_in_port_cell(.PORT_ID_IN(clk_in),
.PORT_ID_OUT(fresh_wire_2));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000020),
.PARAM_PORT_TYPE(2'h0)) config_addr_in_port_cell(.PORT_ID_IN(config_addr_in),
.PORT_ID_OUT(fresh_wire_3));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000020),
.PARAM_PORT_TYPE(2'h0)) config_data_in_port_cell(.PORT_ID_IN(config_data_in),
.PORT_ID_OUT(fresh_wire_4));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) ext_cki_jm_port_cell(.PORT_ID_IN(ext_cki_jm),
.PORT_ID_OUT(fresh_wire_6));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) ext_cki_port_cell(.PORT_ID_IN(ext_cki),
.PORT_ID_OUT(fresh_wire_5));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) ext_ckib_jm_port_cell(.PORT_ID_IN(ext_ckib_jm),
.PORT_ID_OUT(fresh_wire_8));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) ext_ckib_port_cell(.PORT_ID_IN(ext_ckib),
.PORT_ID_OUT(fresh_wire_7));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) ext_frefn_jm_port_cell(.PORT_ID_IN(ext_frefn_jm),
.PORT_ID_OUT(fresh_wire_10));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) ext_frefn_port_cell(.PORT_ID_IN(ext_frefn),
.PORT_ID_OUT(fresh_wire_9));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) ext_frefp_jm_port_cell(.PORT_ID_IN(ext_frefp_jm),
.PORT_ID_OUT(fresh_wire_12));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) ext_frefp_port_cell(.PORT_ID_IN(ext_frefp),
.PORT_ID_OUT(fresh_wire_11));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) ffeed_pad_port_cell(.PORT_ID_IN(fresh_wire_13),
.PORT_ID_OUT(ffeed_pad));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) fout_div_pad_port_cell(.PORT_ID_IN(fresh_wire_14),
.PORT_ID_OUT(fout_div_pad));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) fref_off_pad_port_cell(.PORT_ID_IN(fresh_wire_15),
.PORT_ID_OUT(fref_off_pad));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) frefn_out_jm_port_cell(.PORT_ID_IN(fresh_wire_16),
.PORT_ID_OUT(frefn_out_jm));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) frefp_out_jm_port_cell(.PORT_ID_IN(fresh_wire_17),
.PORT_ID_OUT(frefp_out_jm));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h0000000d),
.PARAM_PORT_TYPE(2'h1)) lf_out_port_cell(.PORT_ID_IN(fresh_wire_18),
.PORT_ID_OUT(lf_out));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(13'h0000),
.PARAM_WIDTH(32'h0000000d)) mdll_top$self_lf_out(.PORT_ID_OUT(fresh_wire_154));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000004),
.PARAM_PORT_TYPE(2'h1)) mdllout_pad_port_cell(.PORT_ID_IN(fresh_wire_19),
.PORT_ID_OUT(mdllout_pad));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$__DOLLAR__and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__memory_core_unq1__DOT__v__COLON__309__DOLLAR__631$op0(.PORT_ID_IN0(fresh_wire_155),
.PORT_ID_IN1(fresh_wire_156),
.PORT_ID_OUT(fresh_wire_157));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$__DOLLAR__and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__memory_core_unq1__DOT__v__COLON__310__DOLLAR__633$op0(.PORT_ID_IN0(fresh_wire_158),
.PORT_ID_IN1(fresh_wire_159),
.PORT_ID_OUT(fresh_wire_160));

	CELL_TYPE_OR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$__DOLLAR__or__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__memory_core_unq1__DOT__v__COLON__309__DOLLAR__630$op0(.PORT_ID_IN0(fresh_wire_161),
.PORT_ID_IN1(fresh_wire_162),
.PORT_ID_OUT(fresh_wire_163));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__471$op0(.PORT_ID_IN0(fresh_wire_164),
.PORT_ID_IN1(fresh_wire_165),
.PORT_ID_OUT(fresh_wire_166));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000002),
.PARAM_OUT_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__206__DOLLAR__488$extendB(.PORT_ID_IN(fresh_wire_167),
.PORT_ID_OUT(fresh_wire_168));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__206__DOLLAR__488$op0(.PORT_ID_IN0(fresh_wire_169),
.PORT_ID_IN1(fresh_wire_170),
.PORT_ID_OUT(fresh_wire_171));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__233__DOLLAR__500$extendA(.PORT_ID_IN(fresh_wire_172),
.PORT_ID_OUT(fresh_wire_173));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__233__DOLLAR__500$op0(.PORT_ID_IN0(fresh_wire_174),
.PORT_ID_IN1(fresh_wire_175),
.PORT_ID_OUT(fresh_wire_176));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__235__DOLLAR__501$extendA(.PORT_ID_IN(fresh_wire_177),
.PORT_ID_OUT(fresh_wire_178));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__235__DOLLAR__501$op0(.PORT_ID_IN0(fresh_wire_179),
.PORT_ID_IN1(fresh_wire_180),
.PORT_ID_OUT(fresh_wire_181));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__242__DOLLAR__504$extendA(.PORT_ID_IN(fresh_wire_182),
.PORT_ID_OUT(fresh_wire_183));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__242__DOLLAR__504$op0(.PORT_ID_IN0(fresh_wire_184),
.PORT_ID_IN1(fresh_wire_185),
.PORT_ID_OUT(fresh_wire_186));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__271__DOLLAR__521$op0(.PORT_ID_IN0(fresh_wire_187),
.PORT_ID_IN1(fresh_wire_188),
.PORT_ID_OUT(fresh_wire_189));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__273__DOLLAR__525$op0(.PORT_ID_IN0(fresh_wire_190),
.PORT_ID_IN1(fresh_wire_191),
.PORT_ID_OUT(fresh_wire_192));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__276__DOLLAR__534$op0(.PORT_ID_IN0(fresh_wire_193),
.PORT_ID_IN1(fresh_wire_194),
.PORT_ID_OUT(fresh_wire_195));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__555$op0(.PORT_ID_IN0(fresh_wire_196),
.PORT_ID_IN1(fresh_wire_197),
.PORT_ID_OUT(fresh_wire_198));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__207__DOLLAR__491$op0(.PORT_ID_IN0(fresh_wire_199),
.PORT_ID_IN1(fresh_wire_200),
.PORT_ID_OUT(fresh_wire_201));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__466$op0(.PORT_ID_IN0(fresh_wire_202),
.PORT_ID_IN1(fresh_wire_203),
.PORT_ID_OUT(fresh_wire_204));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__467$op0(.PORT_ID_IN0(fresh_wire_205),
.PORT_ID_IN1(fresh_wire_206),
.PORT_ID_OUT(fresh_wire_207));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__469$op0(.PORT_ID_IN0(fresh_wire_208),
.PORT_ID_IN1(fresh_wire_209),
.PORT_ID_OUT(fresh_wire_210));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__472$op0(.PORT_ID_IN0(fresh_wire_211),
.PORT_ID_IN1(fresh_wire_212),
.PORT_ID_OUT(fresh_wire_213));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__176__DOLLAR__474$op0(.PORT_ID_IN0(fresh_wire_214),
.PORT_ID_IN1(fresh_wire_215),
.PORT_ID_OUT(fresh_wire_216));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__192__DOLLAR__482$op0(.PORT_ID_IN0(fresh_wire_217),
.PORT_ID_IN1(fresh_wire_218),
.PORT_ID_OUT(fresh_wire_219));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__193__DOLLAR__483$op0(.PORT_ID_IN0(fresh_wire_220),
.PORT_ID_IN1(fresh_wire_221),
.PORT_ID_OUT(fresh_wire_222));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__196__DOLLAR__484$op0(.PORT_ID_IN0(fresh_wire_223),
.PORT_ID_IN1(fresh_wire_224),
.PORT_ID_OUT(fresh_wire_225));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__207__DOLLAR__490$op0(.PORT_ID_IN0(fresh_wire_226),
.PORT_ID_IN1(fresh_wire_227),
.PORT_ID_OUT(fresh_wire_228));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__228__DOLLAR__497$op0(.PORT_ID_IN0(fresh_wire_229),
.PORT_ID_IN1(fresh_wire_230),
.PORT_ID_OUT(fresh_wire_231));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__229__DOLLAR__498$op0(.PORT_ID_IN0(fresh_wire_232),
.PORT_ID_IN1(fresh_wire_233),
.PORT_ID_OUT(fresh_wire_234));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__268__DOLLAR__513$op0(.PORT_ID_IN0(fresh_wire_235),
.PORT_ID_IN1(fresh_wire_236),
.PORT_ID_OUT(fresh_wire_237));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__268__DOLLAR__516$op0(.PORT_ID_IN0(fresh_wire_238),
.PORT_ID_IN1(fresh_wire_239),
.PORT_ID_OUT(fresh_wire_240));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__273__DOLLAR__524$op0(.PORT_ID_IN0(fresh_wire_241),
.PORT_ID_IN1(fresh_wire_242),
.PORT_ID_OUT(fresh_wire_243));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__285__DOLLAR__541$op0(.PORT_ID_IN0(fresh_wire_244),
.PORT_ID_IN1(fresh_wire_245),
.PORT_ID_OUT(fresh_wire_246));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__309__DOLLAR__549$op0(.PORT_ID_IN0(fresh_wire_247),
.PORT_ID_IN1(fresh_wire_248),
.PORT_ID_OUT(fresh_wire_249));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__556$op0(.PORT_ID_IN0(fresh_wire_250),
.PORT_ID_IN1(fresh_wire_251),
.PORT_ID_OUT(fresh_wire_252));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__316__DOLLAR__558$op0(.PORT_ID_IN0(fresh_wire_253),
.PORT_ID_IN1(fresh_wire_254),
.PORT_ID_OUT(fresh_wire_255));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__355__DOLLAR__568$op0(.PORT_ID_IN0(fresh_wire_256),
.PORT_ID_IN1(fresh_wire_257),
.PORT_ID_OUT(fresh_wire_258));

	CELL_TYPE_UGE #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__ge__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__230__DOLLAR__499$op0(.PORT_ID_IN0(fresh_wire_259),
.PORT_ID_IN1(fresh_wire_260),
.PORT_ID_OUT(fresh_wire_261));

	CELL_TYPE_UGE #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__ge__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__239__DOLLAR__503$op0(.PORT_ID_IN0(fresh_wire_262),
.PORT_ID_IN1(fresh_wire_263),
.PORT_ID_OUT(fresh_wire_264));

	CELL_TYPE_UGE #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__ge__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__276__DOLLAR__535$op0(.PORT_ID_IN0(fresh_wire_265),
.PORT_ID_IN1(fresh_wire_266),
.PORT_ID_OUT(fresh_wire_267));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__468$aRed(.PORT_ID_IN(fresh_wire_268),
.PORT_ID_OUT(fresh_wire_269));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__468$andOps(.PORT_ID_IN0(fresh_wire_270),
.PORT_ID_IN1(fresh_wire_271),
.PORT_ID_OUT(fresh_wire_272));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__468$bRed(.PORT_ID_IN(fresh_wire_273),
.PORT_ID_OUT(fresh_wire_274));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__470$aRed(.PORT_ID_IN(fresh_wire_275),
.PORT_ID_OUT(fresh_wire_276));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__470$andOps(.PORT_ID_IN0(fresh_wire_277),
.PORT_ID_IN1(fresh_wire_278),
.PORT_ID_OUT(fresh_wire_279));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__470$bRed(.PORT_ID_IN(fresh_wire_280),
.PORT_ID_OUT(fresh_wire_281));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__473$aRed(.PORT_ID_IN(fresh_wire_282),
.PORT_ID_OUT(fresh_wire_283));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__473$andOps(.PORT_ID_IN0(fresh_wire_284),
.PORT_ID_IN1(fresh_wire_285),
.PORT_ID_OUT(fresh_wire_286));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__473$bRed(.PORT_ID_IN(fresh_wire_287),
.PORT_ID_OUT(fresh_wire_288));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__268__DOLLAR__515$aRed(.PORT_ID_IN(fresh_wire_289),
.PORT_ID_OUT(fresh_wire_290));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__268__DOLLAR__515$andOps(.PORT_ID_IN0(fresh_wire_291),
.PORT_ID_IN1(fresh_wire_292),
.PORT_ID_OUT(fresh_wire_293));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__268__DOLLAR__517$aRed(.PORT_ID_IN(fresh_wire_294),
.PORT_ID_OUT(fresh_wire_295));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__268__DOLLAR__517$andOps(.PORT_ID_IN0(fresh_wire_296),
.PORT_ID_IN1(fresh_wire_297),
.PORT_ID_OUT(fresh_wire_298));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__268__DOLLAR__517$bRed(.PORT_ID_IN(fresh_wire_299),
.PORT_ID_OUT(fresh_wire_300));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__271__DOLLAR__520$aRed(.PORT_ID_IN(fresh_wire_301),
.PORT_ID_OUT(fresh_wire_302));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__271__DOLLAR__520$andOps(.PORT_ID_IN0(fresh_wire_303),
.PORT_ID_IN1(fresh_wire_304),
.PORT_ID_OUT(fresh_wire_305));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__271__DOLLAR__523$aRed(.PORT_ID_IN(fresh_wire_306),
.PORT_ID_OUT(fresh_wire_307));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__271__DOLLAR__523$andOps(.PORT_ID_IN0(fresh_wire_308),
.PORT_ID_IN1(fresh_wire_309),
.PORT_ID_OUT(fresh_wire_310));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__271__DOLLAR__523$bRed(.PORT_ID_IN(fresh_wire_311),
.PORT_ID_OUT(fresh_wire_312));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__276__DOLLAR__536$aRed(.PORT_ID_IN(fresh_wire_313),
.PORT_ID_OUT(fresh_wire_314));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__276__DOLLAR__536$andOps(.PORT_ID_IN0(fresh_wire_315),
.PORT_ID_IN1(fresh_wire_316),
.PORT_ID_OUT(fresh_wire_317));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__276__DOLLAR__536$bRed(.PORT_ID_IN(fresh_wire_318),
.PORT_ID_OUT(fresh_wire_319));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__277__DOLLAR__539$andOps(.PORT_ID_IN0(fresh_wire_320),
.PORT_ID_IN1(fresh_wire_321),
.PORT_ID_OUT(fresh_wire_322));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__277__DOLLAR__539$bRed(.PORT_ID_IN(fresh_wire_323),
.PORT_ID_OUT(fresh_wire_324));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__285__DOLLAR__543$aRed(.PORT_ID_IN(fresh_wire_325),
.PORT_ID_OUT(fresh_wire_326));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__285__DOLLAR__543$andOps(.PORT_ID_IN0(fresh_wire_327),
.PORT_ID_IN1(fresh_wire_328),
.PORT_ID_OUT(fresh_wire_329));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__552$aRed(.PORT_ID_IN(fresh_wire_330),
.PORT_ID_OUT(fresh_wire_331));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__552$andOps(.PORT_ID_IN0(fresh_wire_332),
.PORT_ID_IN1(fresh_wire_333),
.PORT_ID_OUT(fresh_wire_334));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__552$bRed(.PORT_ID_IN(fresh_wire_335),
.PORT_ID_OUT(fresh_wire_336));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__554$aRed(.PORT_ID_IN(fresh_wire_337),
.PORT_ID_OUT(fresh_wire_338));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__554$andOps(.PORT_ID_IN0(fresh_wire_339),
.PORT_ID_IN1(fresh_wire_340),
.PORT_ID_OUT(fresh_wire_341));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__554$bRed(.PORT_ID_IN(fresh_wire_342),
.PORT_ID_OUT(fresh_wire_343));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__557$aRed(.PORT_ID_IN(fresh_wire_344),
.PORT_ID_OUT(fresh_wire_345));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__557$andOps(.PORT_ID_IN0(fresh_wire_346),
.PORT_ID_IN1(fresh_wire_347),
.PORT_ID_OUT(fresh_wire_348));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__557$bRed(.PORT_ID_IN(fresh_wire_349),
.PORT_ID_OUT(fresh_wire_350));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__316__DOLLAR__560$aRed(.PORT_ID_IN(fresh_wire_351),
.PORT_ID_OUT(fresh_wire_352));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__316__DOLLAR__560$andOps(.PORT_ID_IN0(fresh_wire_353),
.PORT_ID_IN1(fresh_wire_354),
.PORT_ID_OUT(fresh_wire_355));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_or__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__344__DOLLAR__565$bRed(.PORT_ID_IN(fresh_wire_356),
.PORT_ID_OUT(fresh_wire_357));

	CELL_TYPE_OR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_or__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__344__DOLLAR__565$orOps(.PORT_ID_IN0(fresh_wire_358),
.PORT_ID_IN1(fresh_wire_359),
.PORT_ID_OUT(fresh_wire_360));

	CELL_TYPE_ULT #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__lt__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__250__DOLLAR__507$op0(.PORT_ID_IN0(fresh_wire_361),
.PORT_ID_IN1(fresh_wire_362),
.PORT_ID_OUT(fresh_wire_363));

	CELL_TYPE_ULT #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__lt__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__271__DOLLAR__522$op0(.PORT_ID_IN0(fresh_wire_364),
.PORT_ID_IN1(fresh_wire_365),
.PORT_ID_OUT(fresh_wire_366));

	CELL_TYPE_NOT #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__not__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__171__DOLLAR__465$op0(.PORT_ID_IN(fresh_wire_367),
.PORT_ID_OUT(fresh_wire_368));

	CELL_TYPE_REG #(.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3712$reg0(.PORT_ID_CLK(fresh_wire_371),
.PORT_ID_IN(fresh_wire_369),
.PORT_ID_OUT(fresh_wire_370));

	CELL_TYPE_REG #(.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(2'hx),
.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3713$reg0(.PORT_ID_CLK(fresh_wire_374),
.PORT_ID_IN(fresh_wire_372),
.PORT_ID_OUT(fresh_wire_373));

	CELL_TYPE_REG #(.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(2'hx),
.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3714$reg0(.PORT_ID_CLK(fresh_wire_377),
.PORT_ID_IN(fresh_wire_375),
.PORT_ID_OUT(fresh_wire_376));

	CELL_TYPE_REG #(.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(16'hxxxx),
.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3716$reg0(.PORT_ID_CLK(fresh_wire_380),
.PORT_ID_IN(fresh_wire_378),
.PORT_ID_OUT(fresh_wire_379));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3718$reg0(.PORT_ID_ARST(fresh_wire_384),
.PORT_ID_CLK(fresh_wire_383),
.PORT_ID_IN(fresh_wire_381),
.PORT_ID_OUT(fresh_wire_382));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3719$reg0(.PORT_ID_ARST(fresh_wire_388),
.PORT_ID_CLK(fresh_wire_387),
.PORT_ID_IN(fresh_wire_385),
.PORT_ID_OUT(fresh_wire_386));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3720$reg0(.PORT_ID_ARST(fresh_wire_392),
.PORT_ID_CLK(fresh_wire_391),
.PORT_ID_IN(fresh_wire_389),
.PORT_ID_OUT(fresh_wire_390));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3721$reg0(.PORT_ID_ARST(fresh_wire_396),
.PORT_ID_CLK(fresh_wire_395),
.PORT_ID_IN(fresh_wire_393),
.PORT_ID_OUT(fresh_wire_394));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3722$reg0(.PORT_ID_ARST(fresh_wire_400),
.PORT_ID_CLK(fresh_wire_399),
.PORT_ID_IN(fresh_wire_397),
.PORT_ID_OUT(fresh_wire_398));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(2'h0),
.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3723$reg0(.PORT_ID_ARST(fresh_wire_404),
.PORT_ID_CLK(fresh_wire_403),
.PORT_ID_IN(fresh_wire_401),
.PORT_ID_OUT(fresh_wire_402));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(16'h0000),
.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3724$reg0(.PORT_ID_ARST(fresh_wire_408),
.PORT_ID_CLK(fresh_wire_407),
.PORT_ID_IN(fresh_wire_405),
.PORT_ID_OUT(fresh_wire_406));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(16'h0000),
.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3725$reg0(.PORT_ID_ARST(fresh_wire_412),
.PORT_ID_CLK(fresh_wire_411),
.PORT_ID_IN(fresh_wire_409),
.PORT_ID_OUT(fresh_wire_410));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(16'h0000),
.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3726$reg0(.PORT_ID_ARST(fresh_wire_416),
.PORT_ID_CLK(fresh_wire_415),
.PORT_ID_IN(fresh_wire_413),
.PORT_ID_OUT(fresh_wire_414));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(16'h0000),
.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3727$reg0(.PORT_ID_ARST(fresh_wire_420),
.PORT_ID_CLK(fresh_wire_419),
.PORT_ID_IN(fresh_wire_417),
.PORT_ID_OUT(fresh_wire_418));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3728$reg0(.PORT_ID_ARST(fresh_wire_424),
.PORT_ID_CLK(fresh_wire_423),
.PORT_ID_IN(fresh_wire_421),
.PORT_ID_OUT(fresh_wire_422));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3729$reg0(.PORT_ID_ARST(fresh_wire_428),
.PORT_ID_CLK(fresh_wire_427),
.PORT_ID_IN(fresh_wire_425),
.PORT_ID_OUT(fresh_wire_426));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3730$reg0(.PORT_ID_ARST(fresh_wire_432),
.PORT_ID_CLK(fresh_wire_431),
.PORT_ID_IN(fresh_wire_429),
.PORT_ID_OUT(fresh_wire_430));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2788$mux0(.PORT_ID_IN0(fresh_wire_433),
.PORT_ID_IN1(fresh_wire_434),
.PORT_ID_OUT(fresh_wire_435),
.PORT_ID_SEL(fresh_wire_436));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2865$mux0(.PORT_ID_IN0(fresh_wire_437),
.PORT_ID_IN1(fresh_wire_438),
.PORT_ID_OUT(fresh_wire_439),
.PORT_ID_SEL(fresh_wire_440));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2867$mux0(.PORT_ID_IN0(fresh_wire_441),
.PORT_ID_IN1(fresh_wire_442),
.PORT_ID_OUT(fresh_wire_443),
.PORT_ID_SEL(fresh_wire_444));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2877$mux0(.PORT_ID_IN0(fresh_wire_445),
.PORT_ID_IN1(fresh_wire_446),
.PORT_ID_OUT(fresh_wire_447),
.PORT_ID_SEL(fresh_wire_448));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2879$mux0(.PORT_ID_IN0(fresh_wire_449),
.PORT_ID_IN1(fresh_wire_450),
.PORT_ID_OUT(fresh_wire_451),
.PORT_ID_SEL(fresh_wire_452));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2888$mux0(.PORT_ID_IN0(fresh_wire_453),
.PORT_ID_IN1(fresh_wire_454),
.PORT_ID_OUT(fresh_wire_455),
.PORT_ID_SEL(fresh_wire_456));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2898$mux0(.PORT_ID_IN0(fresh_wire_457),
.PORT_ID_IN1(fresh_wire_458),
.PORT_ID_OUT(fresh_wire_459),
.PORT_ID_SEL(fresh_wire_460));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2904$mux0(.PORT_ID_IN0(fresh_wire_461),
.PORT_ID_IN1(fresh_wire_462),
.PORT_ID_OUT(fresh_wire_463),
.PORT_ID_SEL(fresh_wire_464));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2907$mux0(.PORT_ID_IN0(fresh_wire_465),
.PORT_ID_IN1(fresh_wire_466),
.PORT_ID_OUT(fresh_wire_467),
.PORT_ID_SEL(fresh_wire_468));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2909$mux0(.PORT_ID_IN0(fresh_wire_469),
.PORT_ID_IN1(fresh_wire_470),
.PORT_ID_OUT(fresh_wire_471),
.PORT_ID_SEL(fresh_wire_472));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2919$mux0(.PORT_ID_IN0(fresh_wire_473),
.PORT_ID_IN1(fresh_wire_474),
.PORT_ID_OUT(fresh_wire_475),
.PORT_ID_SEL(fresh_wire_476));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2923$mux0(.PORT_ID_IN0(fresh_wire_477),
.PORT_ID_IN1(fresh_wire_478),
.PORT_ID_OUT(fresh_wire_479),
.PORT_ID_SEL(fresh_wire_480));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2925$mux0(.PORT_ID_IN0(fresh_wire_481),
.PORT_ID_IN1(fresh_wire_482),
.PORT_ID_OUT(fresh_wire_483),
.PORT_ID_SEL(fresh_wire_484));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2931$mux0(.PORT_ID_IN0(fresh_wire_485),
.PORT_ID_IN1(fresh_wire_486),
.PORT_ID_OUT(fresh_wire_487),
.PORT_ID_SEL(fresh_wire_488));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2934$mux0(.PORT_ID_IN0(fresh_wire_489),
.PORT_ID_IN1(fresh_wire_490),
.PORT_ID_OUT(fresh_wire_491),
.PORT_ID_SEL(fresh_wire_492));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2936$mux0(.PORT_ID_IN0(fresh_wire_493),
.PORT_ID_IN1(fresh_wire_494),
.PORT_ID_OUT(fresh_wire_495),
.PORT_ID_SEL(fresh_wire_496));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2946$mux0(.PORT_ID_IN0(fresh_wire_497),
.PORT_ID_IN1(fresh_wire_498),
.PORT_ID_OUT(fresh_wire_499),
.PORT_ID_SEL(fresh_wire_500));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2952$mux0(.PORT_ID_IN0(fresh_wire_501),
.PORT_ID_IN1(fresh_wire_502),
.PORT_ID_OUT(fresh_wire_503),
.PORT_ID_SEL(fresh_wire_504));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2955$mux0(.PORT_ID_IN0(fresh_wire_505),
.PORT_ID_IN1(fresh_wire_506),
.PORT_ID_OUT(fresh_wire_507),
.PORT_ID_SEL(fresh_wire_508));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2957$mux0(.PORT_ID_IN0(fresh_wire_509),
.PORT_ID_IN1(fresh_wire_510),
.PORT_ID_OUT(fresh_wire_511),
.PORT_ID_SEL(fresh_wire_512));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2967$mux0(.PORT_ID_IN0(fresh_wire_513),
.PORT_ID_IN1(fresh_wire_514),
.PORT_ID_OUT(fresh_wire_515),
.PORT_ID_SEL(fresh_wire_516));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2971$mux0(.PORT_ID_IN0(fresh_wire_517),
.PORT_ID_IN1(fresh_wire_518),
.PORT_ID_OUT(fresh_wire_519),
.PORT_ID_SEL(fresh_wire_520));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2973$mux0(.PORT_ID_IN0(fresh_wire_521),
.PORT_ID_IN1(fresh_wire_522),
.PORT_ID_OUT(fresh_wire_523),
.PORT_ID_SEL(fresh_wire_524));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2979$mux0(.PORT_ID_IN0(fresh_wire_525),
.PORT_ID_IN1(fresh_wire_526),
.PORT_ID_OUT(fresh_wire_527),
.PORT_ID_SEL(fresh_wire_528));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2982$mux0(.PORT_ID_IN0(fresh_wire_529),
.PORT_ID_IN1(fresh_wire_530),
.PORT_ID_OUT(fresh_wire_531),
.PORT_ID_SEL(fresh_wire_532));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2984$mux0(.PORT_ID_IN0(fresh_wire_533),
.PORT_ID_IN1(fresh_wire_534),
.PORT_ID_OUT(fresh_wire_535),
.PORT_ID_SEL(fresh_wire_536));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2993$mux0(.PORT_ID_IN0(fresh_wire_537),
.PORT_ID_IN1(fresh_wire_538),
.PORT_ID_OUT(fresh_wire_539),
.PORT_ID_SEL(fresh_wire_540));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2997$mux0(.PORT_ID_IN0(fresh_wire_541),
.PORT_ID_IN1(fresh_wire_542),
.PORT_ID_OUT(fresh_wire_543),
.PORT_ID_SEL(fresh_wire_544));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2999$mux0(.PORT_ID_IN0(fresh_wire_545),
.PORT_ID_IN1(fresh_wire_546),
.PORT_ID_OUT(fresh_wire_547),
.PORT_ID_SEL(fresh_wire_548));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3013$mux0(.PORT_ID_IN0(fresh_wire_549),
.PORT_ID_IN1(fresh_wire_550),
.PORT_ID_OUT(fresh_wire_551),
.PORT_ID_SEL(fresh_wire_552));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3015$mux0(.PORT_ID_IN0(fresh_wire_553),
.PORT_ID_IN1(fresh_wire_554),
.PORT_ID_OUT(fresh_wire_555),
.PORT_ID_SEL(fresh_wire_556));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3017$mux0(.PORT_ID_IN0(fresh_wire_557),
.PORT_ID_IN1(fresh_wire_558),
.PORT_ID_OUT(fresh_wire_559),
.PORT_ID_SEL(fresh_wire_560));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3033$mux0(.PORT_ID_IN0(fresh_wire_561),
.PORT_ID_IN1(fresh_wire_562),
.PORT_ID_OUT(fresh_wire_563),
.PORT_ID_SEL(fresh_wire_564));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3035$mux0(.PORT_ID_IN0(fresh_wire_565),
.PORT_ID_IN1(fresh_wire_566),
.PORT_ID_OUT(fresh_wire_567),
.PORT_ID_SEL(fresh_wire_568));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3038$mux0(.PORT_ID_IN0(fresh_wire_569),
.PORT_ID_IN1(fresh_wire_570),
.PORT_ID_OUT(fresh_wire_571),
.PORT_ID_SEL(fresh_wire_572));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3057$mux0(.PORT_ID_IN0(fresh_wire_573),
.PORT_ID_IN1(fresh_wire_574),
.PORT_ID_OUT(fresh_wire_575),
.PORT_ID_SEL(fresh_wire_576));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3059$mux0(.PORT_ID_IN0(fresh_wire_577),
.PORT_ID_IN1(fresh_wire_578),
.PORT_ID_OUT(fresh_wire_579),
.PORT_ID_SEL(fresh_wire_580));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3069$mux0(.PORT_ID_IN0(fresh_wire_581),
.PORT_ID_IN1(fresh_wire_582),
.PORT_ID_OUT(fresh_wire_583),
.PORT_ID_SEL(fresh_wire_584));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3072$mux0(.PORT_ID_IN0(fresh_wire_585),
.PORT_ID_IN1(fresh_wire_586),
.PORT_ID_OUT(fresh_wire_587),
.PORT_ID_SEL(fresh_wire_588));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3074$mux0(.PORT_ID_IN0(fresh_wire_589),
.PORT_ID_IN1(fresh_wire_590),
.PORT_ID_OUT(fresh_wire_591),
.PORT_ID_SEL(fresh_wire_592));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__sub__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__244__DOLLAR__505$extendA(.PORT_ID_IN(fresh_wire_593),
.PORT_ID_OUT(fresh_wire_594));

	CELL_TYPE_SUB #(.PARAM_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__sub__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__244__DOLLAR__505$op0(.PORT_ID_IN0(fresh_wire_595),
.PORT_ID_IN1(fresh_wire_596),
.PORT_ID_OUT(fresh_wire_597));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__ternary__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__176__DOLLAR__475$mux0(.PORT_ID_IN0(fresh_wire_598),
.PORT_ID_IN1(fresh_wire_599),
.PORT_ID_OUT(fresh_wire_600),
.PORT_ID_SEL(fresh_wire_601));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__ternary__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__273__DOLLAR__526$mux0(.PORT_ID_IN0(fresh_wire_602),
.PORT_ID_IN1(fresh_wire_603),
.PORT_ID_OUT(fresh_wire_604),
.PORT_ID_SEL(fresh_wire_605));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__ternary__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__273__DOLLAR__526__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(.PORT_ID_OUT(fresh_wire_606));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__ternary__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__355__DOLLAR__569$mux0(.PORT_ID_IN0(fresh_wire_607),
.PORT_ID_IN1(fresh_wire_608),
.PORT_ID_OUT(fresh_wire_609),
.PORT_ID_SEL(fresh_wire_610));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__101__DOLLAR__314$op0(.PORT_ID_IN0(fresh_wire_611),
.PORT_ID_IN1(fresh_wire_612),
.PORT_ID_OUT(fresh_wire_613));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__100__DOLLAR__310$op0(.PORT_ID_IN0(fresh_wire_614),
.PORT_ID_IN1(fresh_wire_615),
.PORT_ID_OUT(fresh_wire_616));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__100__DOLLAR__311$op0(.PORT_ID_IN0(fresh_wire_617),
.PORT_ID_IN1(fresh_wire_618),
.PORT_ID_OUT(fresh_wire_619));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__103__DOLLAR__316$op0(.PORT_ID_IN0(fresh_wire_620),
.PORT_ID_IN1(fresh_wire_621),
.PORT_ID_OUT(fresh_wire_622));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__128__DOLLAR__345$op0(.PORT_ID_IN0(fresh_wire_623),
.PORT_ID_IN1(fresh_wire_624),
.PORT_ID_OUT(fresh_wire_625));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__150__DOLLAR__379$op0(.PORT_ID_IN0(fresh_wire_626),
.PORT_ID_IN1(fresh_wire_627),
.PORT_ID_OUT(fresh_wire_628));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__157__DOLLAR__381$op0(.PORT_ID_IN0(fresh_wire_629),
.PORT_ID_IN1(fresh_wire_630),
.PORT_ID_OUT(fresh_wire_631));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__158__DOLLAR__382$op0(.PORT_ID_IN0(fresh_wire_632),
.PORT_ID_IN1(fresh_wire_633),
.PORT_ID_OUT(fresh_wire_634));

	CELL_TYPE_UGE #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__ge__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__126__DOLLAR__341$op0(.PORT_ID_IN0(fresh_wire_635),
.PORT_ID_IN1(fresh_wire_636),
.PORT_ID_OUT(fresh_wire_637));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__100__DOLLAR__312$aRed(.PORT_ID_IN(fresh_wire_638),
.PORT_ID_OUT(fresh_wire_639));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__100__DOLLAR__312$andOps(.PORT_ID_IN0(fresh_wire_640),
.PORT_ID_IN1(fresh_wire_641),
.PORT_ID_OUT(fresh_wire_642));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__100__DOLLAR__312$bRed(.PORT_ID_IN(fresh_wire_643),
.PORT_ID_OUT(fresh_wire_644));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__100__DOLLAR__313$andOps(.PORT_ID_IN0(fresh_wire_645),
.PORT_ID_IN1(fresh_wire_646),
.PORT_ID_OUT(fresh_wire_647));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__100__DOLLAR__313$bRed(.PORT_ID_IN(fresh_wire_648),
.PORT_ID_OUT(fresh_wire_649));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__103__DOLLAR__317$andOps(.PORT_ID_IN0(fresh_wire_650),
.PORT_ID_IN1(fresh_wire_651),
.PORT_ID_OUT(fresh_wire_652));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__103__DOLLAR__317$bRed(.PORT_ID_IN(fresh_wire_653),
.PORT_ID_OUT(fresh_wire_654));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__125__DOLLAR__340$andOps(.PORT_ID_IN0(fresh_wire_655),
.PORT_ID_IN1(fresh_wire_656),
.PORT_ID_OUT(fresh_wire_657));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__125__DOLLAR__340$bRed(.PORT_ID_IN(fresh_wire_658),
.PORT_ID_OUT(fresh_wire_659));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__127__DOLLAR__344$andOps(.PORT_ID_IN0(fresh_wire_660),
.PORT_ID_IN1(fresh_wire_661),
.PORT_ID_OUT(fresh_wire_662));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__127__DOLLAR__344$bRed(.PORT_ID_IN(fresh_wire_663),
.PORT_ID_OUT(fresh_wire_664));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(2'h0),
.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__procdff__DOLLAR__3739$reg0(.PORT_ID_ARST(fresh_wire_668),
.PORT_ID_CLK(fresh_wire_667),
.PORT_ID_IN(fresh_wire_665),
.PORT_ID_OUT(fresh_wire_666));

	CELL_TYPE_REG #(.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(48'hxxxxxxxxxxxx),
.PARAM_WIDTH(32'h00000030)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__procdff__DOLLAR__3740$reg0(.PORT_ID_CLK(fresh_wire_671),
.PORT_ID_IN(fresh_wire_669),
.PORT_ID_OUT(fresh_wire_670));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3178$mux0(.PORT_ID_IN0(fresh_wire_672),
.PORT_ID_IN1(fresh_wire_673),
.PORT_ID_OUT(fresh_wire_674),
.PORT_ID_SEL(fresh_wire_675));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3181$mux0(.PORT_ID_IN0(fresh_wire_676),
.PORT_ID_IN1(fresh_wire_677),
.PORT_ID_OUT(fresh_wire_678),
.PORT_ID_SEL(fresh_wire_679));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3199$mux0(.PORT_ID_IN0(fresh_wire_680),
.PORT_ID_IN1(fresh_wire_681),
.PORT_ID_OUT(fresh_wire_682),
.PORT_ID_SEL(fresh_wire_683));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3202$mux0(.PORT_ID_IN0(fresh_wire_684),
.PORT_ID_IN1(fresh_wire_685),
.PORT_ID_OUT(fresh_wire_686),
.PORT_ID_SEL(fresh_wire_687));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3211$mux0(.PORT_ID_IN0(fresh_wire_688),
.PORT_ID_IN1(fresh_wire_689),
.PORT_ID_OUT(fresh_wire_690),
.PORT_ID_SEL(fresh_wire_691));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3214$mux0(.PORT_ID_IN0(fresh_wire_692),
.PORT_ID_IN1(fresh_wire_693),
.PORT_ID_OUT(fresh_wire_694),
.PORT_ID_SEL(fresh_wire_695));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3217$mux0(.PORT_ID_IN0(fresh_wire_696),
.PORT_ID_IN1(fresh_wire_697),
.PORT_ID_OUT(fresh_wire_698),
.PORT_ID_SEL(fresh_wire_699));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3219$mux0(.PORT_ID_IN0(fresh_wire_700),
.PORT_ID_IN1(fresh_wire_701),
.PORT_ID_OUT(fresh_wire_702),
.PORT_ID_SEL(fresh_wire_703));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3223$mux0(.PORT_ID_IN0(fresh_wire_704),
.PORT_ID_IN1(fresh_wire_705),
.PORT_ID_OUT(fresh_wire_706),
.PORT_ID_SEL(fresh_wire_707));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3226$mux0(.PORT_ID_IN0(fresh_wire_708),
.PORT_ID_IN1(fresh_wire_709),
.PORT_ID_OUT(fresh_wire_710),
.PORT_ID_SEL(fresh_wire_711));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3228$mux0(.PORT_ID_IN0(fresh_wire_712),
.PORT_ID_IN1(fresh_wire_713),
.PORT_ID_OUT(fresh_wire_714),
.PORT_ID_SEL(fresh_wire_715));

	CELL_TYPE_SUB #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__sub__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__104__DOLLAR__318$op0(.PORT_ID_IN0(fresh_wire_716),
.PORT_ID_IN1(fresh_wire_717),
.PORT_ID_OUT(fresh_wire_718));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__sub__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__110__DOLLAR__326__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(.PORT_ID_OUT(fresh_wire_719));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__103__DOLLAR__747$op0(.PORT_ID_IN0(fresh_wire_720),
.PORT_ID_IN1(fresh_wire_721),
.PORT_ID_OUT(fresh_wire_722));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__106__DOLLAR__751$op0(.PORT_ID_IN0(fresh_wire_723),
.PORT_ID_IN1(fresh_wire_724),
.PORT_ID_OUT(fresh_wire_725));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__102__DOLLAR__744$op0(.PORT_ID_IN0(fresh_wire_726),
.PORT_ID_IN1(fresh_wire_727),
.PORT_ID_OUT(fresh_wire_728));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__102__DOLLAR__745$op0(.PORT_ID_IN0(fresh_wire_729),
.PORT_ID_IN1(fresh_wire_730),
.PORT_ID_OUT(fresh_wire_731));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__105__DOLLAR__748$op0(.PORT_ID_IN0(fresh_wire_732),
.PORT_ID_IN1(fresh_wire_733),
.PORT_ID_OUT(fresh_wire_734));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__108__DOLLAR__753$op0(.PORT_ID_IN0(fresh_wire_735),
.PORT_ID_IN1(fresh_wire_736),
.PORT_ID_OUT(fresh_wire_737));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__120__DOLLAR__760$op0(.PORT_ID_IN0(fresh_wire_738),
.PORT_ID_IN1(fresh_wire_739),
.PORT_ID_OUT(fresh_wire_740));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__120__DOLLAR__761$op0(.PORT_ID_IN0(fresh_wire_741),
.PORT_ID_IN1(fresh_wire_742),
.PORT_ID_OUT(fresh_wire_743));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__133__DOLLAR__784$op0(.PORT_ID_IN0(fresh_wire_744),
.PORT_ID_IN1(fresh_wire_745),
.PORT_ID_OUT(fresh_wire_746));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__135__DOLLAR__785$op0(.PORT_ID_IN0(fresh_wire_747),
.PORT_ID_IN1(fresh_wire_748),
.PORT_ID_OUT(fresh_wire_749));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__137__DOLLAR__786$op0(.PORT_ID_IN0(fresh_wire_750),
.PORT_ID_IN1(fresh_wire_751),
.PORT_ID_OUT(fresh_wire_752));

	CELL_TYPE_UGE #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__ge__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__121__DOLLAR__765$op0(.PORT_ID_IN0(fresh_wire_753),
.PORT_ID_IN1(fresh_wire_754),
.PORT_ID_OUT(fresh_wire_755));

	CELL_TYPE_UGE #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__ge__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__123__DOLLAR__771$op0(.PORT_ID_IN0(fresh_wire_756),
.PORT_ID_IN1(fresh_wire_757),
.PORT_ID_OUT(fresh_wire_758));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__102__DOLLAR__746$aRed(.PORT_ID_IN(fresh_wire_759),
.PORT_ID_OUT(fresh_wire_760));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__102__DOLLAR__746$andOps(.PORT_ID_IN0(fresh_wire_761),
.PORT_ID_IN1(fresh_wire_762),
.PORT_ID_OUT(fresh_wire_763));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__102__DOLLAR__746$bRed(.PORT_ID_IN(fresh_wire_764),
.PORT_ID_OUT(fresh_wire_765));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__105__DOLLAR__750$aRed(.PORT_ID_IN(fresh_wire_766),
.PORT_ID_OUT(fresh_wire_767));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__105__DOLLAR__750$andOps(.PORT_ID_IN0(fresh_wire_768),
.PORT_ID_IN1(fresh_wire_769),
.PORT_ID_OUT(fresh_wire_770));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__105__DOLLAR__750$bRed(.PORT_ID_IN(fresh_wire_771),
.PORT_ID_OUT(fresh_wire_772));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__108__DOLLAR__754$aRed(.PORT_ID_IN(fresh_wire_773),
.PORT_ID_OUT(fresh_wire_774));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__108__DOLLAR__754$andOps(.PORT_ID_IN0(fresh_wire_775),
.PORT_ID_IN1(fresh_wire_776),
.PORT_ID_OUT(fresh_wire_777));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__108__DOLLAR__754$bRed(.PORT_ID_IN(fresh_wire_778),
.PORT_ID_OUT(fresh_wire_779));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__110__DOLLAR__757$aRed(.PORT_ID_IN(fresh_wire_780),
.PORT_ID_OUT(fresh_wire_781));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__110__DOLLAR__757$andOps(.PORT_ID_IN0(fresh_wire_782),
.PORT_ID_IN1(fresh_wire_783),
.PORT_ID_OUT(fresh_wire_784));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__110__DOLLAR__757$bRed(.PORT_ID_IN(fresh_wire_785),
.PORT_ID_OUT(fresh_wire_786));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__120__DOLLAR__762$aRed(.PORT_ID_IN(fresh_wire_787),
.PORT_ID_OUT(fresh_wire_788));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__120__DOLLAR__762$andOps(.PORT_ID_IN0(fresh_wire_789),
.PORT_ID_IN1(fresh_wire_790),
.PORT_ID_OUT(fresh_wire_791));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__120__DOLLAR__762$bRed(.PORT_ID_IN(fresh_wire_792),
.PORT_ID_OUT(fresh_wire_793));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__120__DOLLAR__764$aRed(.PORT_ID_IN(fresh_wire_794),
.PORT_ID_OUT(fresh_wire_795));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__120__DOLLAR__764$andOps(.PORT_ID_IN0(fresh_wire_796),
.PORT_ID_IN1(fresh_wire_797),
.PORT_ID_OUT(fresh_wire_798));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__120__DOLLAR__764$bRed(.PORT_ID_IN(fresh_wire_799),
.PORT_ID_OUT(fresh_wire_800));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__122__DOLLAR__768$aRed(.PORT_ID_IN(fresh_wire_801),
.PORT_ID_OUT(fresh_wire_802));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__122__DOLLAR__768$andOps(.PORT_ID_IN0(fresh_wire_803),
.PORT_ID_IN1(fresh_wire_804),
.PORT_ID_OUT(fresh_wire_805));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__122__DOLLAR__768$bRed(.PORT_ID_IN(fresh_wire_806),
.PORT_ID_OUT(fresh_wire_807));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__122__DOLLAR__770$aRed(.PORT_ID_IN(fresh_wire_808),
.PORT_ID_OUT(fresh_wire_809));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__122__DOLLAR__770$andOps(.PORT_ID_IN0(fresh_wire_810),
.PORT_ID_IN1(fresh_wire_811),
.PORT_ID_OUT(fresh_wire_812));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__122__DOLLAR__770$bRed(.PORT_ID_IN(fresh_wire_813),
.PORT_ID_OUT(fresh_wire_814));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__124__DOLLAR__776$aRed(.PORT_ID_IN(fresh_wire_815),
.PORT_ID_OUT(fresh_wire_816));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__124__DOLLAR__776$andOps(.PORT_ID_IN0(fresh_wire_817),
.PORT_ID_IN1(fresh_wire_818),
.PORT_ID_OUT(fresh_wire_819));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__124__DOLLAR__776$bRed(.PORT_ID_IN(fresh_wire_820),
.PORT_ID_OUT(fresh_wire_821));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__126__DOLLAR__781$aRed(.PORT_ID_IN(fresh_wire_822),
.PORT_ID_OUT(fresh_wire_823));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__126__DOLLAR__781$andOps(.PORT_ID_IN0(fresh_wire_824),
.PORT_ID_IN1(fresh_wire_825),
.PORT_ID_OUT(fresh_wire_826));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__126__DOLLAR__781$bRed(.PORT_ID_IN(fresh_wire_827),
.PORT_ID_OUT(fresh_wire_828));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__99__DOLLAR__740$aRed(.PORT_ID_IN(fresh_wire_829),
.PORT_ID_OUT(fresh_wire_830));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__99__DOLLAR__740$andOps(.PORT_ID_IN0(fresh_wire_831),
.PORT_ID_IN1(fresh_wire_832),
.PORT_ID_OUT(fresh_wire_833));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__99__DOLLAR__740$bRed(.PORT_ID_IN(fresh_wire_834),
.PORT_ID_OUT(fresh_wire_835));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__99__DOLLAR__742$aRed(.PORT_ID_IN(fresh_wire_836),
.PORT_ID_OUT(fresh_wire_837));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__99__DOLLAR__742$andOps(.PORT_ID_IN0(fresh_wire_838),
.PORT_ID_IN1(fresh_wire_839),
.PORT_ID_OUT(fresh_wire_840));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__99__DOLLAR__742$bRed(.PORT_ID_IN(fresh_wire_841),
.PORT_ID_OUT(fresh_wire_842));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_or__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__124__DOLLAR__774$aRed(.PORT_ID_IN(fresh_wire_843),
.PORT_ID_OUT(fresh_wire_844));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_or__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__124__DOLLAR__774$bRed(.PORT_ID_IN(fresh_wire_845),
.PORT_ID_OUT(fresh_wire_846));

	CELL_TYPE_OR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_or__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__124__DOLLAR__774$orOps(.PORT_ID_IN0(fresh_wire_847),
.PORT_ID_IN1(fresh_wire_848),
.PORT_ID_OUT(fresh_wire_849));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_or__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__126__DOLLAR__779$aRed(.PORT_ID_IN(fresh_wire_850),
.PORT_ID_OUT(fresh_wire_851));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_or__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__126__DOLLAR__779$bRed(.PORT_ID_IN(fresh_wire_852),
.PORT_ID_OUT(fresh_wire_853));

	CELL_TYPE_OR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_or__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__126__DOLLAR__779$orOps(.PORT_ID_IN0(fresh_wire_854),
.PORT_ID_IN1(fresh_wire_855),
.PORT_ID_OUT(fresh_wire_856));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(2'h0),
.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procdff__DOLLAR__3701$reg0(.PORT_ID_ARST(fresh_wire_860),
.PORT_ID_CLK(fresh_wire_859),
.PORT_ID_IN(fresh_wire_857),
.PORT_ID_OUT(fresh_wire_858));

	CELL_TYPE_REG #(.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(48'hxxxxxxxxxxxx),
.PARAM_WIDTH(32'h00000030)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procdff__DOLLAR__3702$reg0(.PORT_ID_CLK(fresh_wire_863),
.PORT_ID_IN(fresh_wire_861),
.PORT_ID_OUT(fresh_wire_862));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2382$mux0(.PORT_ID_IN0(fresh_wire_864),
.PORT_ID_IN1(fresh_wire_865),
.PORT_ID_OUT(fresh_wire_866),
.PORT_ID_SEL(fresh_wire_867));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2385$mux0(.PORT_ID_IN0(fresh_wire_868),
.PORT_ID_IN1(fresh_wire_869),
.PORT_ID_OUT(fresh_wire_870),
.PORT_ID_SEL(fresh_wire_871));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2388$mux0(.PORT_ID_IN0(fresh_wire_872),
.PORT_ID_IN1(fresh_wire_873),
.PORT_ID_OUT(fresh_wire_874),
.PORT_ID_SEL(fresh_wire_875));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2390$mux0(.PORT_ID_IN0(fresh_wire_876),
.PORT_ID_IN1(fresh_wire_877),
.PORT_ID_OUT(fresh_wire_878),
.PORT_ID_SEL(fresh_wire_879));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2393$mux0(.PORT_ID_IN0(fresh_wire_880),
.PORT_ID_IN1(fresh_wire_881),
.PORT_ID_OUT(fresh_wire_882),
.PORT_ID_SEL(fresh_wire_883));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2396$mux0(.PORT_ID_IN0(fresh_wire_884),
.PORT_ID_IN1(fresh_wire_885),
.PORT_ID_OUT(fresh_wire_886),
.PORT_ID_SEL(fresh_wire_887));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2399$mux0(.PORT_ID_IN0(fresh_wire_888),
.PORT_ID_IN1(fresh_wire_889),
.PORT_ID_OUT(fresh_wire_890),
.PORT_ID_SEL(fresh_wire_891));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2402$mux0(.PORT_ID_IN0(fresh_wire_892),
.PORT_ID_IN1(fresh_wire_893),
.PORT_ID_OUT(fresh_wire_894),
.PORT_ID_SEL(fresh_wire_895));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2406$mux0(.PORT_ID_IN0(fresh_wire_896),
.PORT_ID_IN1(fresh_wire_897),
.PORT_ID_OUT(fresh_wire_898),
.PORT_ID_SEL(fresh_wire_899));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2409$mux0(.PORT_ID_IN0(fresh_wire_900),
.PORT_ID_IN1(fresh_wire_901),
.PORT_ID_OUT(fresh_wire_902),
.PORT_ID_SEL(fresh_wire_903));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2412$mux0(.PORT_ID_IN0(fresh_wire_904),
.PORT_ID_IN1(fresh_wire_905),
.PORT_ID_OUT(fresh_wire_906),
.PORT_ID_SEL(fresh_wire_907));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2415$mux0(.PORT_ID_IN0(fresh_wire_908),
.PORT_ID_IN1(fresh_wire_909),
.PORT_ID_OUT(fresh_wire_910),
.PORT_ID_SEL(fresh_wire_911));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2418$mux0(.PORT_ID_IN0(fresh_wire_912),
.PORT_ID_IN1(fresh_wire_913),
.PORT_ID_OUT(fresh_wire_914),
.PORT_ID_SEL(fresh_wire_915));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000030)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2427$mux0(.PORT_ID_IN0(fresh_wire_916),
.PORT_ID_IN1(fresh_wire_917),
.PORT_ID_OUT(fresh_wire_918),
.PORT_ID_SEL(fresh_wire_919));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000030)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2430$mux0(.PORT_ID_IN0(fresh_wire_920),
.PORT_ID_IN1(fresh_wire_921),
.PORT_ID_OUT(fresh_wire_922),
.PORT_ID_SEL(fresh_wire_923));

	CELL_TYPE_SUB #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__sub__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__100__DOLLAR__743$op0(.PORT_ID_IN0(fresh_wire_924),
.PORT_ID_IN1(fresh_wire_925),
.PORT_ID_OUT(fresh_wire_926));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__sub__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__100__DOLLAR__743__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(.PORT_ID_OUT(fresh_wire_927));

	CELL_TYPE_NOT #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$__DOLLAR__not__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__mem_unq1__DOT__v__COLON__65__DOLLAR__575$op0(.PORT_ID_IN(fresh_wire_928),
.PORT_ID_OUT(fresh_wire_929));

	CELL_TYPE_NOT #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$__DOLLAR__not__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__mem_unq1__DOT__v__COLON__66__DOLLAR__576$op0(.PORT_ID_IN(fresh_wire_930),
.PORT_ID_OUT(fresh_wire_931));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__sram_512w_16b__DOT__v__COLON__38__DOLLAR__1114$op0(.PORT_ID_IN0(fresh_wire_932),
.PORT_ID_IN1(fresh_wire_933),
.PORT_ID_OUT(fresh_wire_934));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__sram_512w_16b__DOT__v__COLON__40__DOLLAR__1116$op0(.PORT_ID_IN0(fresh_wire_935),
.PORT_ID_IN1(fresh_wire_936),
.PORT_ID_OUT(fresh_wire_937));

	CELL_TYPE_REG #(.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(16'hxxxx),
.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procdff__DOLLAR__3630$reg0(.PORT_ID_CLK(fresh_wire_940),
.PORT_ID_IN(fresh_wire_938),
.PORT_ID_OUT(fresh_wire_939));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1557$mux0(.PORT_ID_IN0(fresh_wire_941),
.PORT_ID_IN1(fresh_wire_942),
.PORT_ID_OUT(fresh_wire_943),
.PORT_ID_SEL(fresh_wire_944));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1567$mux0(.PORT_ID_IN0(fresh_wire_945),
.PORT_ID_IN1(fresh_wire_946),
.PORT_ID_OUT(fresh_wire_947),
.PORT_ID_SEL(fresh_wire_948));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1567__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(.PORT_ID_OUT(fresh_wire_949));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1569$mux0(.PORT_ID_IN0(fresh_wire_950),
.PORT_ID_IN1(fresh_wire_951),
.PORT_ID_OUT(fresh_wire_952),
.PORT_ID_SEL(fresh_wire_953));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576$mux0(.PORT_ID_IN0(fresh_wire_954),
.PORT_ID_IN1(fresh_wire_955),
.PORT_ID_OUT(fresh_wire_956),
.PORT_ID_SEL(fresh_wire_957));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0$uConst(.PORT_ID_OUT(fresh_wire_958));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10$uConst(.PORT_ID_OUT(fresh_wire_959));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11$uConst(.PORT_ID_OUT(fresh_wire_960));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12$uConst(.PORT_ID_OUT(fresh_wire_961));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13$uConst(.PORT_ID_OUT(fresh_wire_962));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14$uConst(.PORT_ID_OUT(fresh_wire_963));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15$uConst(.PORT_ID_OUT(fresh_wire_964));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1$uConst(.PORT_ID_OUT(fresh_wire_965));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2$uConst(.PORT_ID_OUT(fresh_wire_966));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3$uConst(.PORT_ID_OUT(fresh_wire_967));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4$uConst(.PORT_ID_OUT(fresh_wire_968));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5$uConst(.PORT_ID_OUT(fresh_wire_969));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6$uConst(.PORT_ID_OUT(fresh_wire_970));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7$uConst(.PORT_ID_OUT(fresh_wire_971));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8$uConst(.PORT_ID_OUT(fresh_wire_972));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9$uConst(.PORT_ID_OUT(fresh_wire_973));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578$mux0(.PORT_ID_IN0(fresh_wire_974),
.PORT_ID_IN1(fresh_wire_975),
.PORT_ID_OUT(fresh_wire_976),
.PORT_ID_SEL(fresh_wire_977));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0$uConst(.PORT_ID_OUT(fresh_wire_978));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10$uConst(.PORT_ID_OUT(fresh_wire_979));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11$uConst(.PORT_ID_OUT(fresh_wire_980));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12$uConst(.PORT_ID_OUT(fresh_wire_981));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13$uConst(.PORT_ID_OUT(fresh_wire_982));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14$uConst(.PORT_ID_OUT(fresh_wire_983));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15$uConst(.PORT_ID_OUT(fresh_wire_984));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1$uConst(.PORT_ID_OUT(fresh_wire_985));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2$uConst(.PORT_ID_OUT(fresh_wire_986));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3$uConst(.PORT_ID_OUT(fresh_wire_987));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4$uConst(.PORT_ID_OUT(fresh_wire_988));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5$uConst(.PORT_ID_OUT(fresh_wire_989));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6$uConst(.PORT_ID_OUT(fresh_wire_990));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7$uConst(.PORT_ID_OUT(fresh_wire_991));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8$uConst(.PORT_ID_OUT(fresh_wire_992));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9$uConst(.PORT_ID_OUT(fresh_wire_993));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000009)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585$mux0(.PORT_ID_IN0(fresh_wire_994),
.PORT_ID_IN1(fresh_wire_995),
.PORT_ID_OUT(fresh_wire_996),
.PORT_ID_SEL(fresh_wire_997));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0$uConst(.PORT_ID_OUT(fresh_wire_998));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1$uConst(.PORT_ID_OUT(fresh_wire_999));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2$uConst(.PORT_ID_OUT(fresh_wire_1000));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3$uConst(.PORT_ID_OUT(fresh_wire_1001));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4$uConst(.PORT_ID_OUT(fresh_wire_1002));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5$uConst(.PORT_ID_OUT(fresh_wire_1003));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6$uConst(.PORT_ID_OUT(fresh_wire_1004));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7$uConst(.PORT_ID_OUT(fresh_wire_1005));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8$uConst(.PORT_ID_OUT(fresh_wire_1006));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000009)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587$mux0(.PORT_ID_IN0(fresh_wire_1007),
.PORT_ID_IN1(fresh_wire_1008),
.PORT_ID_OUT(fresh_wire_1009),
.PORT_ID_SEL(fresh_wire_1010));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0$uConst(.PORT_ID_OUT(fresh_wire_1011));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1$uConst(.PORT_ID_OUT(fresh_wire_1012));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2$uConst(.PORT_ID_OUT(fresh_wire_1013));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3$uConst(.PORT_ID_OUT(fresh_wire_1014));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4$uConst(.PORT_ID_OUT(fresh_wire_1015));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5$uConst(.PORT_ID_OUT(fresh_wire_1016));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6$uConst(.PORT_ID_OUT(fresh_wire_1017));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7$uConst(.PORT_ID_OUT(fresh_wire_1018));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8$uConst(.PORT_ID_OUT(fresh_wire_1019));

	CELL_TYPE_MEM #(.PARAM_HAS_INIT(1'h0),
.PARAM_MEM_DEPTH(32'h00000200),
.PARAM_MEM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst0$mem_inst$data_array$mem(.PORT_ID_CLK(fresh_wire_1020),
.PORT_ID_RADDR(fresh_wire_1021),
.PORT_ID_RDATA(fresh_wire_1022),
.PORT_ID_WADDR(fresh_wire_1023),
.PORT_ID_WDATA(fresh_wire_1024),
.PORT_ID_WEN(fresh_wire_1025));

	CELL_TYPE_NOT #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$__DOLLAR__not__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__mem_unq1__DOT__v__COLON__65__DOLLAR__575$op0(.PORT_ID_IN(fresh_wire_1026),
.PORT_ID_OUT(fresh_wire_1027));

	CELL_TYPE_NOT #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$__DOLLAR__not__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__mem_unq1__DOT__v__COLON__66__DOLLAR__576$op0(.PORT_ID_IN(fresh_wire_1028),
.PORT_ID_OUT(fresh_wire_1029));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__sram_512w_16b__DOT__v__COLON__38__DOLLAR__1114$op0(.PORT_ID_IN0(fresh_wire_1030),
.PORT_ID_IN1(fresh_wire_1031),
.PORT_ID_OUT(fresh_wire_1032));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__sram_512w_16b__DOT__v__COLON__40__DOLLAR__1116$op0(.PORT_ID_IN0(fresh_wire_1033),
.PORT_ID_IN1(fresh_wire_1034),
.PORT_ID_OUT(fresh_wire_1035));

	CELL_TYPE_REG #(.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(16'hxxxx),
.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procdff__DOLLAR__3630$reg0(.PORT_ID_CLK(fresh_wire_1038),
.PORT_ID_IN(fresh_wire_1036),
.PORT_ID_OUT(fresh_wire_1037));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1557$mux0(.PORT_ID_IN0(fresh_wire_1039),
.PORT_ID_IN1(fresh_wire_1040),
.PORT_ID_OUT(fresh_wire_1041),
.PORT_ID_SEL(fresh_wire_1042));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1567$mux0(.PORT_ID_IN0(fresh_wire_1043),
.PORT_ID_IN1(fresh_wire_1044),
.PORT_ID_OUT(fresh_wire_1045),
.PORT_ID_SEL(fresh_wire_1046));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1567__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(.PORT_ID_OUT(fresh_wire_1047));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1569$mux0(.PORT_ID_IN0(fresh_wire_1048),
.PORT_ID_IN1(fresh_wire_1049),
.PORT_ID_OUT(fresh_wire_1050),
.PORT_ID_SEL(fresh_wire_1051));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576$mux0(.PORT_ID_IN0(fresh_wire_1052),
.PORT_ID_IN1(fresh_wire_1053),
.PORT_ID_OUT(fresh_wire_1054),
.PORT_ID_SEL(fresh_wire_1055));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0$uConst(.PORT_ID_OUT(fresh_wire_1056));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10$uConst(.PORT_ID_OUT(fresh_wire_1057));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11$uConst(.PORT_ID_OUT(fresh_wire_1058));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12$uConst(.PORT_ID_OUT(fresh_wire_1059));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13$uConst(.PORT_ID_OUT(fresh_wire_1060));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14$uConst(.PORT_ID_OUT(fresh_wire_1061));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15$uConst(.PORT_ID_OUT(fresh_wire_1062));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1$uConst(.PORT_ID_OUT(fresh_wire_1063));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2$uConst(.PORT_ID_OUT(fresh_wire_1064));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3$uConst(.PORT_ID_OUT(fresh_wire_1065));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4$uConst(.PORT_ID_OUT(fresh_wire_1066));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5$uConst(.PORT_ID_OUT(fresh_wire_1067));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6$uConst(.PORT_ID_OUT(fresh_wire_1068));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7$uConst(.PORT_ID_OUT(fresh_wire_1069));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8$uConst(.PORT_ID_OUT(fresh_wire_1070));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9$uConst(.PORT_ID_OUT(fresh_wire_1071));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578$mux0(.PORT_ID_IN0(fresh_wire_1072),
.PORT_ID_IN1(fresh_wire_1073),
.PORT_ID_OUT(fresh_wire_1074),
.PORT_ID_SEL(fresh_wire_1075));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0$uConst(.PORT_ID_OUT(fresh_wire_1076));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10$uConst(.PORT_ID_OUT(fresh_wire_1077));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11$uConst(.PORT_ID_OUT(fresh_wire_1078));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12$uConst(.PORT_ID_OUT(fresh_wire_1079));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13$uConst(.PORT_ID_OUT(fresh_wire_1080));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14$uConst(.PORT_ID_OUT(fresh_wire_1081));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15$uConst(.PORT_ID_OUT(fresh_wire_1082));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1$uConst(.PORT_ID_OUT(fresh_wire_1083));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2$uConst(.PORT_ID_OUT(fresh_wire_1084));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3$uConst(.PORT_ID_OUT(fresh_wire_1085));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4$uConst(.PORT_ID_OUT(fresh_wire_1086));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5$uConst(.PORT_ID_OUT(fresh_wire_1087));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6$uConst(.PORT_ID_OUT(fresh_wire_1088));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7$uConst(.PORT_ID_OUT(fresh_wire_1089));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8$uConst(.PORT_ID_OUT(fresh_wire_1090));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9$uConst(.PORT_ID_OUT(fresh_wire_1091));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000009)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585$mux0(.PORT_ID_IN0(fresh_wire_1092),
.PORT_ID_IN1(fresh_wire_1093),
.PORT_ID_OUT(fresh_wire_1094),
.PORT_ID_SEL(fresh_wire_1095));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0$uConst(.PORT_ID_OUT(fresh_wire_1096));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1$uConst(.PORT_ID_OUT(fresh_wire_1097));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2$uConst(.PORT_ID_OUT(fresh_wire_1098));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3$uConst(.PORT_ID_OUT(fresh_wire_1099));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4$uConst(.PORT_ID_OUT(fresh_wire_1100));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5$uConst(.PORT_ID_OUT(fresh_wire_1101));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6$uConst(.PORT_ID_OUT(fresh_wire_1102));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7$uConst(.PORT_ID_OUT(fresh_wire_1103));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8$uConst(.PORT_ID_OUT(fresh_wire_1104));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000009)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587$mux0(.PORT_ID_IN0(fresh_wire_1105),
.PORT_ID_IN1(fresh_wire_1106),
.PORT_ID_OUT(fresh_wire_1107),
.PORT_ID_SEL(fresh_wire_1108));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0$uConst(.PORT_ID_OUT(fresh_wire_1109));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1$uConst(.PORT_ID_OUT(fresh_wire_1110));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2$uConst(.PORT_ID_OUT(fresh_wire_1111));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3$uConst(.PORT_ID_OUT(fresh_wire_1112));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4$uConst(.PORT_ID_OUT(fresh_wire_1113));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5$uConst(.PORT_ID_OUT(fresh_wire_1114));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6$uConst(.PORT_ID_OUT(fresh_wire_1115));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7$uConst(.PORT_ID_OUT(fresh_wire_1116));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8$uConst(.PORT_ID_OUT(fresh_wire_1117));

	CELL_TYPE_MEM #(.PARAM_HAS_INIT(1'h0),
.PARAM_MEM_DEPTH(32'h00000200),
.PARAM_MEM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst1$mem_inst$data_array$mem(.PORT_ID_CLK(fresh_wire_1118),
.PORT_ID_RADDR(fresh_wire_1119),
.PORT_ID_RDATA(fresh_wire_1120),
.PORT_ID_WADDR(fresh_wire_1121),
.PORT_ID_WDATA(fresh_wire_1122),
.PORT_ID_WEN(fresh_wire_1123));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T0_in_port_cell(.PORT_ID_IN(pad_S0_T0_in),
.PORT_ID_OUT(fresh_wire_20));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T0_out_port_cell(.PORT_ID_IN(fresh_wire_21),
.PORT_ID_OUT(pad_S0_T0_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T10_in_port_cell(.PORT_ID_IN(pad_S0_T10_in),
.PORT_ID_OUT(fresh_wire_22));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T10_out_port_cell(.PORT_ID_IN(fresh_wire_23),
.PORT_ID_OUT(pad_S0_T10_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T11_in_port_cell(.PORT_ID_IN(pad_S0_T11_in),
.PORT_ID_OUT(fresh_wire_24));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T11_out_port_cell(.PORT_ID_IN(fresh_wire_25),
.PORT_ID_OUT(pad_S0_T11_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T12_in_port_cell(.PORT_ID_IN(pad_S0_T12_in),
.PORT_ID_OUT(fresh_wire_26));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T12_out_port_cell(.PORT_ID_IN(fresh_wire_27),
.PORT_ID_OUT(pad_S0_T12_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T13_in_port_cell(.PORT_ID_IN(pad_S0_T13_in),
.PORT_ID_OUT(fresh_wire_28));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T13_out_port_cell(.PORT_ID_IN(fresh_wire_29),
.PORT_ID_OUT(pad_S0_T13_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T14_in_port_cell(.PORT_ID_IN(pad_S0_T14_in),
.PORT_ID_OUT(fresh_wire_30));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T14_out_port_cell(.PORT_ID_IN(fresh_wire_31),
.PORT_ID_OUT(pad_S0_T14_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T15_in_port_cell(.PORT_ID_IN(pad_S0_T15_in),
.PORT_ID_OUT(fresh_wire_32));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T15_out_port_cell(.PORT_ID_IN(fresh_wire_33),
.PORT_ID_OUT(pad_S0_T15_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T1_in_port_cell(.PORT_ID_IN(pad_S0_T1_in),
.PORT_ID_OUT(fresh_wire_34));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T1_out_port_cell(.PORT_ID_IN(fresh_wire_35),
.PORT_ID_OUT(pad_S0_T1_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T2_in_port_cell(.PORT_ID_IN(pad_S0_T2_in),
.PORT_ID_OUT(fresh_wire_36));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T2_out_port_cell(.PORT_ID_IN(fresh_wire_37),
.PORT_ID_OUT(pad_S0_T2_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T3_in_port_cell(.PORT_ID_IN(pad_S0_T3_in),
.PORT_ID_OUT(fresh_wire_38));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T3_out_port_cell(.PORT_ID_IN(fresh_wire_39),
.PORT_ID_OUT(pad_S0_T3_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T4_in_port_cell(.PORT_ID_IN(pad_S0_T4_in),
.PORT_ID_OUT(fresh_wire_40));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T4_out_port_cell(.PORT_ID_IN(fresh_wire_41),
.PORT_ID_OUT(pad_S0_T4_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T5_in_port_cell(.PORT_ID_IN(pad_S0_T5_in),
.PORT_ID_OUT(fresh_wire_42));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T5_out_port_cell(.PORT_ID_IN(fresh_wire_43),
.PORT_ID_OUT(pad_S0_T5_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T6_in_port_cell(.PORT_ID_IN(pad_S0_T6_in),
.PORT_ID_OUT(fresh_wire_44));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T6_out_port_cell(.PORT_ID_IN(fresh_wire_45),
.PORT_ID_OUT(pad_S0_T6_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T7_in_port_cell(.PORT_ID_IN(pad_S0_T7_in),
.PORT_ID_OUT(fresh_wire_46));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T7_out_port_cell(.PORT_ID_IN(fresh_wire_47),
.PORT_ID_OUT(pad_S0_T7_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T8_in_port_cell(.PORT_ID_IN(pad_S0_T8_in),
.PORT_ID_OUT(fresh_wire_48));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T8_out_port_cell(.PORT_ID_IN(fresh_wire_49),
.PORT_ID_OUT(pad_S0_T8_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T9_in_port_cell(.PORT_ID_IN(pad_S0_T9_in),
.PORT_ID_OUT(fresh_wire_50));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T9_out_port_cell(.PORT_ID_IN(fresh_wire_51),
.PORT_ID_OUT(pad_S0_T9_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T0_in_port_cell(.PORT_ID_IN(pad_S1_T0_in),
.PORT_ID_OUT(fresh_wire_52));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T0_out_port_cell(.PORT_ID_IN(fresh_wire_53),
.PORT_ID_OUT(pad_S1_T0_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T10_in_port_cell(.PORT_ID_IN(pad_S1_T10_in),
.PORT_ID_OUT(fresh_wire_54));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T10_out_port_cell(.PORT_ID_IN(fresh_wire_55),
.PORT_ID_OUT(pad_S1_T10_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T11_in_port_cell(.PORT_ID_IN(pad_S1_T11_in),
.PORT_ID_OUT(fresh_wire_56));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T11_out_port_cell(.PORT_ID_IN(fresh_wire_57),
.PORT_ID_OUT(pad_S1_T11_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T12_in_port_cell(.PORT_ID_IN(pad_S1_T12_in),
.PORT_ID_OUT(fresh_wire_58));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T12_out_port_cell(.PORT_ID_IN(fresh_wire_59),
.PORT_ID_OUT(pad_S1_T12_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T13_in_port_cell(.PORT_ID_IN(pad_S1_T13_in),
.PORT_ID_OUT(fresh_wire_60));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T13_out_port_cell(.PORT_ID_IN(fresh_wire_61),
.PORT_ID_OUT(pad_S1_T13_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T14_in_port_cell(.PORT_ID_IN(pad_S1_T14_in),
.PORT_ID_OUT(fresh_wire_62));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T14_out_port_cell(.PORT_ID_IN(fresh_wire_63),
.PORT_ID_OUT(pad_S1_T14_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T15_in_port_cell(.PORT_ID_IN(pad_S1_T15_in),
.PORT_ID_OUT(fresh_wire_64));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T15_out_port_cell(.PORT_ID_IN(fresh_wire_65),
.PORT_ID_OUT(pad_S1_T15_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T1_in_port_cell(.PORT_ID_IN(pad_S1_T1_in),
.PORT_ID_OUT(fresh_wire_66));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T1_out_port_cell(.PORT_ID_IN(fresh_wire_67),
.PORT_ID_OUT(pad_S1_T1_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T2_in_port_cell(.PORT_ID_IN(pad_S1_T2_in),
.PORT_ID_OUT(fresh_wire_68));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T2_out_port_cell(.PORT_ID_IN(fresh_wire_69),
.PORT_ID_OUT(pad_S1_T2_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T3_in_port_cell(.PORT_ID_IN(pad_S1_T3_in),
.PORT_ID_OUT(fresh_wire_70));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T3_out_port_cell(.PORT_ID_IN(fresh_wire_71),
.PORT_ID_OUT(pad_S1_T3_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T4_in_port_cell(.PORT_ID_IN(pad_S1_T4_in),
.PORT_ID_OUT(fresh_wire_72));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T4_out_port_cell(.PORT_ID_IN(fresh_wire_73),
.PORT_ID_OUT(pad_S1_T4_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T5_in_port_cell(.PORT_ID_IN(pad_S1_T5_in),
.PORT_ID_OUT(fresh_wire_74));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T5_out_port_cell(.PORT_ID_IN(fresh_wire_75),
.PORT_ID_OUT(pad_S1_T5_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T6_in_port_cell(.PORT_ID_IN(pad_S1_T6_in),
.PORT_ID_OUT(fresh_wire_76));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T6_out_port_cell(.PORT_ID_IN(fresh_wire_77),
.PORT_ID_OUT(pad_S1_T6_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T7_in_port_cell(.PORT_ID_IN(pad_S1_T7_in),
.PORT_ID_OUT(fresh_wire_78));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T7_out_port_cell(.PORT_ID_IN(fresh_wire_79),
.PORT_ID_OUT(pad_S1_T7_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T8_in_port_cell(.PORT_ID_IN(pad_S1_T8_in),
.PORT_ID_OUT(fresh_wire_80));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T8_out_port_cell(.PORT_ID_IN(fresh_wire_81),
.PORT_ID_OUT(pad_S1_T8_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T9_in_port_cell(.PORT_ID_IN(pad_S1_T9_in),
.PORT_ID_OUT(fresh_wire_82));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T9_out_port_cell(.PORT_ID_IN(fresh_wire_83),
.PORT_ID_OUT(pad_S1_T9_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T0_in_port_cell(.PORT_ID_IN(pad_S2_T0_in),
.PORT_ID_OUT(fresh_wire_84));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T0_out_port_cell(.PORT_ID_IN(fresh_wire_85),
.PORT_ID_OUT(pad_S2_T0_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T10_in_port_cell(.PORT_ID_IN(pad_S2_T10_in),
.PORT_ID_OUT(fresh_wire_86));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T10_out_port_cell(.PORT_ID_IN(fresh_wire_87),
.PORT_ID_OUT(pad_S2_T10_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T11_in_port_cell(.PORT_ID_IN(pad_S2_T11_in),
.PORT_ID_OUT(fresh_wire_88));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T11_out_port_cell(.PORT_ID_IN(fresh_wire_89),
.PORT_ID_OUT(pad_S2_T11_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T12_in_port_cell(.PORT_ID_IN(pad_S2_T12_in),
.PORT_ID_OUT(fresh_wire_90));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T12_out_port_cell(.PORT_ID_IN(fresh_wire_91),
.PORT_ID_OUT(pad_S2_T12_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T13_in_port_cell(.PORT_ID_IN(pad_S2_T13_in),
.PORT_ID_OUT(fresh_wire_92));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T13_out_port_cell(.PORT_ID_IN(fresh_wire_93),
.PORT_ID_OUT(pad_S2_T13_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T14_in_port_cell(.PORT_ID_IN(pad_S2_T14_in),
.PORT_ID_OUT(fresh_wire_94));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T14_out_port_cell(.PORT_ID_IN(fresh_wire_95),
.PORT_ID_OUT(pad_S2_T14_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T15_in_port_cell(.PORT_ID_IN(pad_S2_T15_in),
.PORT_ID_OUT(fresh_wire_96));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T15_out_port_cell(.PORT_ID_IN(fresh_wire_97),
.PORT_ID_OUT(pad_S2_T15_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T1_in_port_cell(.PORT_ID_IN(pad_S2_T1_in),
.PORT_ID_OUT(fresh_wire_98));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T1_out_port_cell(.PORT_ID_IN(fresh_wire_99),
.PORT_ID_OUT(pad_S2_T1_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T2_in_port_cell(.PORT_ID_IN(pad_S2_T2_in),
.PORT_ID_OUT(fresh_wire_100));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T2_out_port_cell(.PORT_ID_IN(fresh_wire_101),
.PORT_ID_OUT(pad_S2_T2_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T3_in_port_cell(.PORT_ID_IN(pad_S2_T3_in),
.PORT_ID_OUT(fresh_wire_102));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T3_out_port_cell(.PORT_ID_IN(fresh_wire_103),
.PORT_ID_OUT(pad_S2_T3_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T4_in_port_cell(.PORT_ID_IN(pad_S2_T4_in),
.PORT_ID_OUT(fresh_wire_104));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T4_out_port_cell(.PORT_ID_IN(fresh_wire_105),
.PORT_ID_OUT(pad_S2_T4_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T5_in_port_cell(.PORT_ID_IN(pad_S2_T5_in),
.PORT_ID_OUT(fresh_wire_106));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T5_out_port_cell(.PORT_ID_IN(fresh_wire_107),
.PORT_ID_OUT(pad_S2_T5_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T6_in_port_cell(.PORT_ID_IN(pad_S2_T6_in),
.PORT_ID_OUT(fresh_wire_108));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T6_out_port_cell(.PORT_ID_IN(fresh_wire_109),
.PORT_ID_OUT(pad_S2_T6_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T7_in_port_cell(.PORT_ID_IN(pad_S2_T7_in),
.PORT_ID_OUT(fresh_wire_110));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T7_out_port_cell(.PORT_ID_IN(fresh_wire_111),
.PORT_ID_OUT(pad_S2_T7_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T8_in_port_cell(.PORT_ID_IN(pad_S2_T8_in),
.PORT_ID_OUT(fresh_wire_112));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T8_out_port_cell(.PORT_ID_IN(fresh_wire_113),
.PORT_ID_OUT(pad_S2_T8_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T9_in_port_cell(.PORT_ID_IN(pad_S2_T9_in),
.PORT_ID_OUT(fresh_wire_114));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T9_out_port_cell(.PORT_ID_IN(fresh_wire_115),
.PORT_ID_OUT(pad_S2_T9_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T0_in_port_cell(.PORT_ID_IN(pad_S3_T0_in),
.PORT_ID_OUT(fresh_wire_116));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T0_out_port_cell(.PORT_ID_IN(fresh_wire_117),
.PORT_ID_OUT(pad_S3_T0_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T10_in_port_cell(.PORT_ID_IN(pad_S3_T10_in),
.PORT_ID_OUT(fresh_wire_118));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T10_out_port_cell(.PORT_ID_IN(fresh_wire_119),
.PORT_ID_OUT(pad_S3_T10_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T11_in_port_cell(.PORT_ID_IN(pad_S3_T11_in),
.PORT_ID_OUT(fresh_wire_120));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T11_out_port_cell(.PORT_ID_IN(fresh_wire_121),
.PORT_ID_OUT(pad_S3_T11_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T12_in_port_cell(.PORT_ID_IN(pad_S3_T12_in),
.PORT_ID_OUT(fresh_wire_122));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T12_out_port_cell(.PORT_ID_IN(fresh_wire_123),
.PORT_ID_OUT(pad_S3_T12_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T13_in_port_cell(.PORT_ID_IN(pad_S3_T13_in),
.PORT_ID_OUT(fresh_wire_124));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T13_out_port_cell(.PORT_ID_IN(fresh_wire_125),
.PORT_ID_OUT(pad_S3_T13_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T14_in_port_cell(.PORT_ID_IN(pad_S3_T14_in),
.PORT_ID_OUT(fresh_wire_126));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T14_out_port_cell(.PORT_ID_IN(fresh_wire_127),
.PORT_ID_OUT(pad_S3_T14_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T15_in_port_cell(.PORT_ID_IN(pad_S3_T15_in),
.PORT_ID_OUT(fresh_wire_128));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T15_out_port_cell(.PORT_ID_IN(fresh_wire_129),
.PORT_ID_OUT(pad_S3_T15_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T1_in_port_cell(.PORT_ID_IN(pad_S3_T1_in),
.PORT_ID_OUT(fresh_wire_130));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T1_out_port_cell(.PORT_ID_IN(fresh_wire_131),
.PORT_ID_OUT(pad_S3_T1_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T2_in_port_cell(.PORT_ID_IN(pad_S3_T2_in),
.PORT_ID_OUT(fresh_wire_132));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T2_out_port_cell(.PORT_ID_IN(fresh_wire_133),
.PORT_ID_OUT(pad_S3_T2_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T3_in_port_cell(.PORT_ID_IN(pad_S3_T3_in),
.PORT_ID_OUT(fresh_wire_134));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T3_out_port_cell(.PORT_ID_IN(fresh_wire_135),
.PORT_ID_OUT(pad_S3_T3_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T4_in_port_cell(.PORT_ID_IN(pad_S3_T4_in),
.PORT_ID_OUT(fresh_wire_136));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T4_out_port_cell(.PORT_ID_IN(fresh_wire_137),
.PORT_ID_OUT(pad_S3_T4_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T5_in_port_cell(.PORT_ID_IN(pad_S3_T5_in),
.PORT_ID_OUT(fresh_wire_138));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T5_out_port_cell(.PORT_ID_IN(fresh_wire_139),
.PORT_ID_OUT(pad_S3_T5_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T6_in_port_cell(.PORT_ID_IN(pad_S3_T6_in),
.PORT_ID_OUT(fresh_wire_140));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T6_out_port_cell(.PORT_ID_IN(fresh_wire_141),
.PORT_ID_OUT(pad_S3_T6_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T7_in_port_cell(.PORT_ID_IN(pad_S3_T7_in),
.PORT_ID_OUT(fresh_wire_142));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T7_out_port_cell(.PORT_ID_IN(fresh_wire_143),
.PORT_ID_OUT(pad_S3_T7_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T8_in_port_cell(.PORT_ID_IN(pad_S3_T8_in),
.PORT_ID_OUT(fresh_wire_144));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T8_out_port_cell(.PORT_ID_IN(fresh_wire_145),
.PORT_ID_OUT(pad_S3_T8_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T9_in_port_cell(.PORT_ID_IN(pad_S3_T9_in),
.PORT_ID_OUT(fresh_wire_146));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T9_out_port_cell(.PORT_ID_IN(fresh_wire_147),
.PORT_ID_OUT(pad_S3_T9_out));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000011),
.PARAM_OUT_WIDTH(32'h00000022)) pe_0x15$test_pe$test_pe_comp$test_mult_add$__DOLLAR__mul__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__1503$extendA(.PORT_ID_IN(fresh_wire_1124),
.PORT_ID_OUT(fresh_wire_1125));

	CELL_TYPE_MUL #(.PARAM_WIDTH(32'h00000022)) pe_0x15$test_pe$test_pe_comp$test_mult_add$__DOLLAR__mul__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__1503$op0(.PORT_ID_IN0(fresh_wire_1126),
.PORT_ID_IN1(fresh_wire_1127),
.PORT_ID_OUT(fresh_wire_1128));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000011)) pe_0x16$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$extendA(.PORT_ID_IN(fresh_wire_1129),
.PORT_ID_OUT(fresh_wire_1130));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000011)) pe_0x16$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$op0(.PORT_ID_IN0(fresh_wire_1131),
.PORT_ID_IN1(fresh_wire_1132),
.PORT_ID_OUT(fresh_wire_1133));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000011)) pe_0x16$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1495$op0(.PORT_ID_IN0(fresh_wire_1134),
.PORT_ID_IN1(fresh_wire_1135),
.PORT_ID_OUT(fresh_wire_1136));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000011),
.PARAM_OUT_WIDTH(32'h00000022)) pe_0x17$test_pe$test_pe_comp$test_mult_add$__DOLLAR__mul__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__1503$extendA(.PORT_ID_IN(fresh_wire_1137),
.PORT_ID_OUT(fresh_wire_1138));

	CELL_TYPE_MUL #(.PARAM_WIDTH(32'h00000022)) pe_0x17$test_pe$test_pe_comp$test_mult_add$__DOLLAR__mul__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__1503$op0(.PORT_ID_IN0(fresh_wire_1139),
.PORT_ID_IN1(fresh_wire_1140),
.PORT_ID_OUT(fresh_wire_1141));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000011)) pe_0x29$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$extendA(.PORT_ID_IN(fresh_wire_1142),
.PORT_ID_OUT(fresh_wire_1143));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000011)) pe_0x29$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$extendB(.PORT_ID_IN(fresh_wire_1144),
.PORT_ID_OUT(fresh_wire_1145));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000011)) pe_0x29$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$op0(.PORT_ID_IN0(fresh_wire_1146),
.PORT_ID_IN1(fresh_wire_1147),
.PORT_ID_OUT(fresh_wire_1148));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000011)) pe_0x29$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1495$op0(.PORT_ID_IN0(fresh_wire_1149),
.PORT_ID_IN1(fresh_wire_1150),
.PORT_ID_OUT(fresh_wire_1151));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) pe_0xFF__DOT__tile_id__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(.PORT_ID_OUT(fresh_wire_1152));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) reset_in_port_cell(.PORT_ID_IN(reset_in),
.PORT_ID_OUT(fresh_wire_148));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) tck_port_cell(.PORT_ID_IN(tck),
.PORT_ID_OUT(fresh_wire_149));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) tdi_port_cell(.PORT_ID_IN(tdi),
.PORT_ID_OUT(fresh_wire_150));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) tdo_port_cell(.PORT_ID_IN(fresh_wire_151),
.PORT_ID_OUT(tdo));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) tms_port_cell(.PORT_ID_IN(tms),
.PORT_ID_OUT(fresh_wire_152));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) trst_n_port_cell(.PORT_ID_IN(trst_n),
.PORT_ID_OUT(fresh_wire_153));

	assign fresh_wire_0[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_13[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_14[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_15[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_16[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_17[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_18[ 0 ] = fresh_wire_154[ 0 ];
	assign fresh_wire_18[ 1 ] = fresh_wire_154[ 1 ];
	assign fresh_wire_18[ 2 ] = fresh_wire_154[ 2 ];
	assign fresh_wire_18[ 3 ] = fresh_wire_154[ 3 ];
	assign fresh_wire_18[ 4 ] = fresh_wire_154[ 4 ];
	assign fresh_wire_18[ 5 ] = fresh_wire_154[ 5 ];
	assign fresh_wire_18[ 6 ] = fresh_wire_154[ 6 ];
	assign fresh_wire_18[ 7 ] = fresh_wire_154[ 7 ];
	assign fresh_wire_18[ 8 ] = fresh_wire_154[ 8 ];
	assign fresh_wire_18[ 9 ] = fresh_wire_154[ 9 ];
	assign fresh_wire_18[ 10 ] = fresh_wire_154[ 10 ];
	assign fresh_wire_18[ 11 ] = fresh_wire_154[ 11 ];
	assign fresh_wire_18[ 12 ] = fresh_wire_154[ 12 ];
	assign fresh_wire_19[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_19[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_19[ 2 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_19[ 3 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_21[ 0 ] = fresh_wire_1151[ 15 ];
	assign fresh_wire_23[ 0 ] = fresh_wire_1151[ 5 ];
	assign fresh_wire_25[ 0 ] = fresh_wire_1151[ 4 ];
	assign fresh_wire_27[ 0 ] = fresh_wire_1151[ 3 ];
	assign fresh_wire_29[ 0 ] = fresh_wire_1151[ 2 ];
	assign fresh_wire_31[ 0 ] = fresh_wire_1151[ 1 ];
	assign fresh_wire_33[ 0 ] = fresh_wire_1151[ 0 ];
	assign fresh_wire_35[ 0 ] = fresh_wire_1151[ 14 ];
	assign fresh_wire_37[ 0 ] = fresh_wire_1151[ 13 ];
	assign fresh_wire_39[ 0 ] = fresh_wire_1151[ 12 ];
	assign fresh_wire_41[ 0 ] = fresh_wire_1151[ 11 ];
	assign fresh_wire_43[ 0 ] = fresh_wire_1151[ 10 ];
	assign fresh_wire_45[ 0 ] = fresh_wire_1151[ 9 ];
	assign fresh_wire_47[ 0 ] = fresh_wire_1151[ 8 ];
	assign fresh_wire_49[ 0 ] = fresh_wire_1151[ 7 ];
	assign fresh_wire_51[ 0 ] = fresh_wire_1151[ 6 ];
	assign fresh_wire_53[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_55[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_57[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_59[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_61[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_63[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_65[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_67[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_69[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_71[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_73[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_75[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_77[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_79[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_81[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_83[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_85[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_87[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_89[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_91[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_93[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_95[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_97[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_99[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_101[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_103[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_105[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_107[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_109[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_111[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_113[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_115[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_117[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_119[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_121[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_123[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_125[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_127[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_129[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_131[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_133[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_135[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_137[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_139[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_141[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_143[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_145[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_147[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_151[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_155[ 0 ] = fresh_wire_1169[ 0 ];
	assign fresh_wire_156[ 0 ] = fresh_wire_163[ 0 ];
	assign fresh_wire_158[ 0 ] = fresh_wire_1169[ 0 ];
	assign fresh_wire_159[ 0 ] = fresh_wire_163[ 0 ];
	assign fresh_wire_161[ 0 ] = fresh_wire_426[ 0 ];
	assign fresh_wire_162[ 0 ] = fresh_wire_201[ 0 ];
	assign fresh_wire_164[ 0 ] = fresh_wire_406[ 0 ];
	assign fresh_wire_164[ 1 ] = fresh_wire_406[ 1 ];
	assign fresh_wire_164[ 2 ] = fresh_wire_406[ 2 ];
	assign fresh_wire_164[ 3 ] = fresh_wire_406[ 3 ];
	assign fresh_wire_164[ 4 ] = fresh_wire_406[ 4 ];
	assign fresh_wire_164[ 5 ] = fresh_wire_406[ 5 ];
	assign fresh_wire_164[ 6 ] = fresh_wire_406[ 6 ];
	assign fresh_wire_164[ 7 ] = fresh_wire_406[ 7 ];
	assign fresh_wire_164[ 8 ] = fresh_wire_406[ 8 ];
	assign fresh_wire_164[ 9 ] = fresh_wire_406[ 9 ];
	assign fresh_wire_164[ 10 ] = fresh_wire_406[ 10 ];
	assign fresh_wire_164[ 11 ] = fresh_wire_406[ 11 ];
	assign fresh_wire_164[ 12 ] = fresh_wire_406[ 12 ];
	assign fresh_wire_164[ 13 ] = fresh_wire_406[ 13 ];
	assign fresh_wire_164[ 14 ] = fresh_wire_406[ 14 ];
	assign fresh_wire_164[ 15 ] = fresh_wire_406[ 15 ];
	assign fresh_wire_165[ 0 ] = fresh_wire_1154[ 0 ];
	assign fresh_wire_165[ 1 ] = fresh_wire_1154[ 1 ];
	assign fresh_wire_165[ 2 ] = fresh_wire_1154[ 2 ];
	assign fresh_wire_165[ 3 ] = fresh_wire_1154[ 3 ];
	assign fresh_wire_165[ 4 ] = fresh_wire_1154[ 4 ];
	assign fresh_wire_165[ 5 ] = fresh_wire_1154[ 5 ];
	assign fresh_wire_165[ 6 ] = fresh_wire_1154[ 6 ];
	assign fresh_wire_165[ 7 ] = fresh_wire_1154[ 7 ];
	assign fresh_wire_165[ 8 ] = fresh_wire_1154[ 8 ];
	assign fresh_wire_165[ 9 ] = fresh_wire_1154[ 9 ];
	assign fresh_wire_165[ 10 ] = fresh_wire_1154[ 10 ];
	assign fresh_wire_165[ 11 ] = fresh_wire_1154[ 11 ];
	assign fresh_wire_165[ 12 ] = fresh_wire_1154[ 12 ];
	assign fresh_wire_165[ 13 ] = fresh_wire_1154[ 13 ];
	assign fresh_wire_165[ 14 ] = fresh_wire_1154[ 14 ];
	assign fresh_wire_165[ 15 ] = fresh_wire_1154[ 15 ];
	assign fresh_wire_167[ 0 ] = fresh_wire_666[ 0 ];
	assign fresh_wire_167[ 1 ] = fresh_wire_666[ 1 ];
	assign fresh_wire_169[ 0 ] = fresh_wire_418[ 0 ];
	assign fresh_wire_169[ 1 ] = fresh_wire_418[ 1 ];
	assign fresh_wire_169[ 2 ] = fresh_wire_418[ 2 ];
	assign fresh_wire_169[ 3 ] = fresh_wire_418[ 3 ];
	assign fresh_wire_169[ 4 ] = fresh_wire_418[ 4 ];
	assign fresh_wire_169[ 5 ] = fresh_wire_418[ 5 ];
	assign fresh_wire_169[ 6 ] = fresh_wire_418[ 6 ];
	assign fresh_wire_169[ 7 ] = fresh_wire_418[ 7 ];
	assign fresh_wire_169[ 8 ] = fresh_wire_418[ 8 ];
	assign fresh_wire_169[ 9 ] = fresh_wire_418[ 9 ];
	assign fresh_wire_169[ 10 ] = fresh_wire_418[ 10 ];
	assign fresh_wire_169[ 11 ] = fresh_wire_418[ 11 ];
	assign fresh_wire_169[ 12 ] = fresh_wire_418[ 12 ];
	assign fresh_wire_169[ 13 ] = fresh_wire_418[ 13 ];
	assign fresh_wire_169[ 14 ] = fresh_wire_418[ 14 ];
	assign fresh_wire_169[ 15 ] = fresh_wire_418[ 15 ];
	assign fresh_wire_170[ 0 ] = fresh_wire_168[ 0 ];
	assign fresh_wire_170[ 1 ] = fresh_wire_168[ 1 ];
	assign fresh_wire_170[ 2 ] = fresh_wire_168[ 2 ];
	assign fresh_wire_170[ 3 ] = fresh_wire_168[ 3 ];
	assign fresh_wire_170[ 4 ] = fresh_wire_168[ 4 ];
	assign fresh_wire_170[ 5 ] = fresh_wire_168[ 5 ];
	assign fresh_wire_170[ 6 ] = fresh_wire_168[ 6 ];
	assign fresh_wire_170[ 7 ] = fresh_wire_168[ 7 ];
	assign fresh_wire_170[ 8 ] = fresh_wire_168[ 8 ];
	assign fresh_wire_170[ 9 ] = fresh_wire_168[ 9 ];
	assign fresh_wire_170[ 10 ] = fresh_wire_168[ 10 ];
	assign fresh_wire_170[ 11 ] = fresh_wire_168[ 11 ];
	assign fresh_wire_170[ 12 ] = fresh_wire_168[ 12 ];
	assign fresh_wire_170[ 13 ] = fresh_wire_168[ 13 ];
	assign fresh_wire_170[ 14 ] = fresh_wire_168[ 14 ];
	assign fresh_wire_170[ 15 ] = fresh_wire_168[ 15 ];
	assign fresh_wire_172[ 0 ] = fresh_wire_414[ 0 ];
	assign fresh_wire_172[ 1 ] = fresh_wire_414[ 1 ];
	assign fresh_wire_172[ 2 ] = fresh_wire_414[ 2 ];
	assign fresh_wire_172[ 3 ] = fresh_wire_414[ 3 ];
	assign fresh_wire_172[ 4 ] = fresh_wire_414[ 4 ];
	assign fresh_wire_172[ 5 ] = fresh_wire_414[ 5 ];
	assign fresh_wire_172[ 6 ] = fresh_wire_414[ 6 ];
	assign fresh_wire_172[ 7 ] = fresh_wire_414[ 7 ];
	assign fresh_wire_172[ 8 ] = fresh_wire_414[ 8 ];
	assign fresh_wire_172[ 9 ] = fresh_wire_414[ 9 ];
	assign fresh_wire_172[ 10 ] = fresh_wire_414[ 10 ];
	assign fresh_wire_172[ 11 ] = fresh_wire_414[ 11 ];
	assign fresh_wire_172[ 12 ] = fresh_wire_414[ 12 ];
	assign fresh_wire_172[ 13 ] = fresh_wire_414[ 13 ];
	assign fresh_wire_172[ 14 ] = fresh_wire_414[ 14 ];
	assign fresh_wire_172[ 15 ] = fresh_wire_414[ 15 ];
	assign fresh_wire_174[ 0 ] = fresh_wire_173[ 0 ];
	assign fresh_wire_174[ 1 ] = fresh_wire_173[ 1 ];
	assign fresh_wire_174[ 2 ] = fresh_wire_173[ 2 ];
	assign fresh_wire_174[ 3 ] = fresh_wire_173[ 3 ];
	assign fresh_wire_174[ 4 ] = fresh_wire_173[ 4 ];
	assign fresh_wire_174[ 5 ] = fresh_wire_173[ 5 ];
	assign fresh_wire_174[ 6 ] = fresh_wire_173[ 6 ];
	assign fresh_wire_174[ 7 ] = fresh_wire_173[ 7 ];
	assign fresh_wire_174[ 8 ] = fresh_wire_173[ 8 ];
	assign fresh_wire_174[ 9 ] = fresh_wire_173[ 9 ];
	assign fresh_wire_174[ 10 ] = fresh_wire_173[ 10 ];
	assign fresh_wire_174[ 11 ] = fresh_wire_173[ 11 ];
	assign fresh_wire_174[ 12 ] = fresh_wire_173[ 12 ];
	assign fresh_wire_174[ 13 ] = fresh_wire_173[ 13 ];
	assign fresh_wire_174[ 14 ] = fresh_wire_173[ 14 ];
	assign fresh_wire_174[ 15 ] = fresh_wire_173[ 15 ];
	assign fresh_wire_174[ 16 ] = fresh_wire_173[ 16 ];
	assign fresh_wire_174[ 17 ] = fresh_wire_173[ 17 ];
	assign fresh_wire_174[ 18 ] = fresh_wire_173[ 18 ];
	assign fresh_wire_174[ 19 ] = fresh_wire_173[ 19 ];
	assign fresh_wire_174[ 20 ] = fresh_wire_173[ 20 ];
	assign fresh_wire_174[ 21 ] = fresh_wire_173[ 21 ];
	assign fresh_wire_174[ 22 ] = fresh_wire_173[ 22 ];
	assign fresh_wire_174[ 23 ] = fresh_wire_173[ 23 ];
	assign fresh_wire_174[ 24 ] = fresh_wire_173[ 24 ];
	assign fresh_wire_174[ 25 ] = fresh_wire_173[ 25 ];
	assign fresh_wire_174[ 26 ] = fresh_wire_173[ 26 ];
	assign fresh_wire_174[ 27 ] = fresh_wire_173[ 27 ];
	assign fresh_wire_174[ 28 ] = fresh_wire_173[ 28 ];
	assign fresh_wire_174[ 29 ] = fresh_wire_173[ 29 ];
	assign fresh_wire_174[ 30 ] = fresh_wire_173[ 30 ];
	assign fresh_wire_174[ 31 ] = fresh_wire_173[ 31 ];
	assign fresh_wire_175[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_175[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 2 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 3 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 4 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 5 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 6 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 7 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 8 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 9 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 10 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 11 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 12 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 13 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 14 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 15 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 16 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 17 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 18 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 19 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 20 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 21 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 22 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 23 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 24 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 25 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 26 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 27 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 28 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 29 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 30 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_175[ 31 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_177[ 0 ] = fresh_wire_418[ 0 ];
	assign fresh_wire_177[ 1 ] = fresh_wire_418[ 1 ];
	assign fresh_wire_177[ 2 ] = fresh_wire_418[ 2 ];
	assign fresh_wire_177[ 3 ] = fresh_wire_418[ 3 ];
	assign fresh_wire_177[ 4 ] = fresh_wire_418[ 4 ];
	assign fresh_wire_177[ 5 ] = fresh_wire_418[ 5 ];
	assign fresh_wire_177[ 6 ] = fresh_wire_418[ 6 ];
	assign fresh_wire_177[ 7 ] = fresh_wire_418[ 7 ];
	assign fresh_wire_177[ 8 ] = fresh_wire_418[ 8 ];
	assign fresh_wire_177[ 9 ] = fresh_wire_418[ 9 ];
	assign fresh_wire_177[ 10 ] = fresh_wire_418[ 10 ];
	assign fresh_wire_177[ 11 ] = fresh_wire_418[ 11 ];
	assign fresh_wire_177[ 12 ] = fresh_wire_418[ 12 ];
	assign fresh_wire_177[ 13 ] = fresh_wire_418[ 13 ];
	assign fresh_wire_177[ 14 ] = fresh_wire_418[ 14 ];
	assign fresh_wire_177[ 15 ] = fresh_wire_418[ 15 ];
	assign fresh_wire_179[ 0 ] = fresh_wire_178[ 0 ];
	assign fresh_wire_179[ 1 ] = fresh_wire_178[ 1 ];
	assign fresh_wire_179[ 2 ] = fresh_wire_178[ 2 ];
	assign fresh_wire_179[ 3 ] = fresh_wire_178[ 3 ];
	assign fresh_wire_179[ 4 ] = fresh_wire_178[ 4 ];
	assign fresh_wire_179[ 5 ] = fresh_wire_178[ 5 ];
	assign fresh_wire_179[ 6 ] = fresh_wire_178[ 6 ];
	assign fresh_wire_179[ 7 ] = fresh_wire_178[ 7 ];
	assign fresh_wire_179[ 8 ] = fresh_wire_178[ 8 ];
	assign fresh_wire_179[ 9 ] = fresh_wire_178[ 9 ];
	assign fresh_wire_179[ 10 ] = fresh_wire_178[ 10 ];
	assign fresh_wire_179[ 11 ] = fresh_wire_178[ 11 ];
	assign fresh_wire_179[ 12 ] = fresh_wire_178[ 12 ];
	assign fresh_wire_179[ 13 ] = fresh_wire_178[ 13 ];
	assign fresh_wire_179[ 14 ] = fresh_wire_178[ 14 ];
	assign fresh_wire_179[ 15 ] = fresh_wire_178[ 15 ];
	assign fresh_wire_179[ 16 ] = fresh_wire_178[ 16 ];
	assign fresh_wire_179[ 17 ] = fresh_wire_178[ 17 ];
	assign fresh_wire_179[ 18 ] = fresh_wire_178[ 18 ];
	assign fresh_wire_179[ 19 ] = fresh_wire_178[ 19 ];
	assign fresh_wire_179[ 20 ] = fresh_wire_178[ 20 ];
	assign fresh_wire_179[ 21 ] = fresh_wire_178[ 21 ];
	assign fresh_wire_179[ 22 ] = fresh_wire_178[ 22 ];
	assign fresh_wire_179[ 23 ] = fresh_wire_178[ 23 ];
	assign fresh_wire_179[ 24 ] = fresh_wire_178[ 24 ];
	assign fresh_wire_179[ 25 ] = fresh_wire_178[ 25 ];
	assign fresh_wire_179[ 26 ] = fresh_wire_178[ 26 ];
	assign fresh_wire_179[ 27 ] = fresh_wire_178[ 27 ];
	assign fresh_wire_179[ 28 ] = fresh_wire_178[ 28 ];
	assign fresh_wire_179[ 29 ] = fresh_wire_178[ 29 ];
	assign fresh_wire_179[ 30 ] = fresh_wire_178[ 30 ];
	assign fresh_wire_179[ 31 ] = fresh_wire_178[ 31 ];
	assign fresh_wire_180[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 1 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_180[ 2 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 3 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 4 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 5 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 6 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 7 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 8 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 9 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 10 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 11 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 12 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 13 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 14 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 15 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 16 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 17 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 18 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 19 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 20 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 21 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 22 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 23 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 24 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 25 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 26 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 27 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 28 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 29 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 30 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_180[ 31 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_182[ 0 ] = fresh_wire_410[ 0 ];
	assign fresh_wire_182[ 1 ] = fresh_wire_410[ 1 ];
	assign fresh_wire_182[ 2 ] = fresh_wire_410[ 2 ];
	assign fresh_wire_182[ 3 ] = fresh_wire_410[ 3 ];
	assign fresh_wire_182[ 4 ] = fresh_wire_410[ 4 ];
	assign fresh_wire_182[ 5 ] = fresh_wire_410[ 5 ];
	assign fresh_wire_182[ 6 ] = fresh_wire_410[ 6 ];
	assign fresh_wire_182[ 7 ] = fresh_wire_410[ 7 ];
	assign fresh_wire_182[ 8 ] = fresh_wire_410[ 8 ];
	assign fresh_wire_182[ 9 ] = fresh_wire_410[ 9 ];
	assign fresh_wire_182[ 10 ] = fresh_wire_410[ 10 ];
	assign fresh_wire_182[ 11 ] = fresh_wire_410[ 11 ];
	assign fresh_wire_182[ 12 ] = fresh_wire_410[ 12 ];
	assign fresh_wire_182[ 13 ] = fresh_wire_410[ 13 ];
	assign fresh_wire_182[ 14 ] = fresh_wire_410[ 14 ];
	assign fresh_wire_182[ 15 ] = fresh_wire_410[ 15 ];
	assign fresh_wire_184[ 0 ] = fresh_wire_183[ 0 ];
	assign fresh_wire_184[ 1 ] = fresh_wire_183[ 1 ];
	assign fresh_wire_184[ 2 ] = fresh_wire_183[ 2 ];
	assign fresh_wire_184[ 3 ] = fresh_wire_183[ 3 ];
	assign fresh_wire_184[ 4 ] = fresh_wire_183[ 4 ];
	assign fresh_wire_184[ 5 ] = fresh_wire_183[ 5 ];
	assign fresh_wire_184[ 6 ] = fresh_wire_183[ 6 ];
	assign fresh_wire_184[ 7 ] = fresh_wire_183[ 7 ];
	assign fresh_wire_184[ 8 ] = fresh_wire_183[ 8 ];
	assign fresh_wire_184[ 9 ] = fresh_wire_183[ 9 ];
	assign fresh_wire_184[ 10 ] = fresh_wire_183[ 10 ];
	assign fresh_wire_184[ 11 ] = fresh_wire_183[ 11 ];
	assign fresh_wire_184[ 12 ] = fresh_wire_183[ 12 ];
	assign fresh_wire_184[ 13 ] = fresh_wire_183[ 13 ];
	assign fresh_wire_184[ 14 ] = fresh_wire_183[ 14 ];
	assign fresh_wire_184[ 15 ] = fresh_wire_183[ 15 ];
	assign fresh_wire_184[ 16 ] = fresh_wire_183[ 16 ];
	assign fresh_wire_184[ 17 ] = fresh_wire_183[ 17 ];
	assign fresh_wire_184[ 18 ] = fresh_wire_183[ 18 ];
	assign fresh_wire_184[ 19 ] = fresh_wire_183[ 19 ];
	assign fresh_wire_184[ 20 ] = fresh_wire_183[ 20 ];
	assign fresh_wire_184[ 21 ] = fresh_wire_183[ 21 ];
	assign fresh_wire_184[ 22 ] = fresh_wire_183[ 22 ];
	assign fresh_wire_184[ 23 ] = fresh_wire_183[ 23 ];
	assign fresh_wire_184[ 24 ] = fresh_wire_183[ 24 ];
	assign fresh_wire_184[ 25 ] = fresh_wire_183[ 25 ];
	assign fresh_wire_184[ 26 ] = fresh_wire_183[ 26 ];
	assign fresh_wire_184[ 27 ] = fresh_wire_183[ 27 ];
	assign fresh_wire_184[ 28 ] = fresh_wire_183[ 28 ];
	assign fresh_wire_184[ 29 ] = fresh_wire_183[ 29 ];
	assign fresh_wire_184[ 30 ] = fresh_wire_183[ 30 ];
	assign fresh_wire_184[ 31 ] = fresh_wire_183[ 31 ];
	assign fresh_wire_185[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_185[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 2 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 3 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 4 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 5 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 6 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 7 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 8 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 9 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 10 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 11 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 12 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 13 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 14 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 15 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 16 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 17 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 18 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 19 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 20 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 21 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 22 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 23 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 24 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 25 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 26 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 27 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 28 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 29 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 30 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_185[ 31 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_187[ 0 ] = fresh_wire_406[ 0 ];
	assign fresh_wire_187[ 1 ] = fresh_wire_406[ 1 ];
	assign fresh_wire_187[ 2 ] = fresh_wire_406[ 2 ];
	assign fresh_wire_187[ 3 ] = fresh_wire_406[ 3 ];
	assign fresh_wire_187[ 4 ] = fresh_wire_406[ 4 ];
	assign fresh_wire_187[ 5 ] = fresh_wire_406[ 5 ];
	assign fresh_wire_187[ 6 ] = fresh_wire_406[ 6 ];
	assign fresh_wire_187[ 7 ] = fresh_wire_406[ 7 ];
	assign fresh_wire_187[ 8 ] = fresh_wire_406[ 8 ];
	assign fresh_wire_187[ 9 ] = fresh_wire_406[ 9 ];
	assign fresh_wire_187[ 10 ] = fresh_wire_406[ 10 ];
	assign fresh_wire_187[ 11 ] = fresh_wire_406[ 11 ];
	assign fresh_wire_187[ 12 ] = fresh_wire_406[ 12 ];
	assign fresh_wire_187[ 13 ] = fresh_wire_406[ 13 ];
	assign fresh_wire_187[ 14 ] = fresh_wire_406[ 14 ];
	assign fresh_wire_187[ 15 ] = fresh_wire_406[ 15 ];
	assign fresh_wire_188[ 0 ] = fresh_wire_1155[ 0 ];
	assign fresh_wire_188[ 1 ] = fresh_wire_1155[ 1 ];
	assign fresh_wire_188[ 2 ] = fresh_wire_1155[ 2 ];
	assign fresh_wire_188[ 3 ] = fresh_wire_1155[ 3 ];
	assign fresh_wire_188[ 4 ] = fresh_wire_1155[ 4 ];
	assign fresh_wire_188[ 5 ] = fresh_wire_1155[ 5 ];
	assign fresh_wire_188[ 6 ] = fresh_wire_1155[ 6 ];
	assign fresh_wire_188[ 7 ] = fresh_wire_1155[ 7 ];
	assign fresh_wire_188[ 8 ] = fresh_wire_1155[ 8 ];
	assign fresh_wire_188[ 9 ] = fresh_wire_1155[ 9 ];
	assign fresh_wire_188[ 10 ] = fresh_wire_1155[ 10 ];
	assign fresh_wire_188[ 11 ] = fresh_wire_1155[ 11 ];
	assign fresh_wire_188[ 12 ] = fresh_wire_1155[ 12 ];
	assign fresh_wire_188[ 13 ] = fresh_wire_1155[ 13 ];
	assign fresh_wire_188[ 14 ] = fresh_wire_1155[ 14 ];
	assign fresh_wire_188[ 15 ] = fresh_wire_1155[ 15 ];
	assign fresh_wire_190[ 0 ] = fresh_wire_406[ 0 ];
	assign fresh_wire_190[ 1 ] = fresh_wire_406[ 1 ];
	assign fresh_wire_190[ 2 ] = fresh_wire_406[ 2 ];
	assign fresh_wire_190[ 3 ] = fresh_wire_406[ 3 ];
	assign fresh_wire_190[ 4 ] = fresh_wire_406[ 4 ];
	assign fresh_wire_190[ 5 ] = fresh_wire_406[ 5 ];
	assign fresh_wire_190[ 6 ] = fresh_wire_406[ 6 ];
	assign fresh_wire_190[ 7 ] = fresh_wire_406[ 7 ];
	assign fresh_wire_190[ 8 ] = fresh_wire_406[ 8 ];
	assign fresh_wire_190[ 9 ] = fresh_wire_406[ 9 ];
	assign fresh_wire_190[ 10 ] = fresh_wire_406[ 10 ];
	assign fresh_wire_190[ 11 ] = fresh_wire_406[ 11 ];
	assign fresh_wire_190[ 12 ] = fresh_wire_406[ 12 ];
	assign fresh_wire_190[ 13 ] = fresh_wire_406[ 13 ];
	assign fresh_wire_190[ 14 ] = fresh_wire_406[ 14 ];
	assign fresh_wire_190[ 15 ] = fresh_wire_406[ 15 ];
	assign fresh_wire_191[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_191[ 1 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_191[ 2 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_191[ 3 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_191[ 4 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_191[ 5 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_191[ 6 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_191[ 7 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_191[ 8 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_191[ 9 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_191[ 10 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_191[ 11 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_191[ 12 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_191[ 13 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_191[ 14 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_191[ 15 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_193[ 0 ] = fresh_wire_406[ 0 ];
	assign fresh_wire_193[ 1 ] = fresh_wire_406[ 1 ];
	assign fresh_wire_193[ 2 ] = fresh_wire_406[ 2 ];
	assign fresh_wire_193[ 3 ] = fresh_wire_406[ 3 ];
	assign fresh_wire_193[ 4 ] = fresh_wire_406[ 4 ];
	assign fresh_wire_193[ 5 ] = fresh_wire_406[ 5 ];
	assign fresh_wire_193[ 6 ] = fresh_wire_406[ 6 ];
	assign fresh_wire_193[ 7 ] = fresh_wire_406[ 7 ];
	assign fresh_wire_193[ 8 ] = fresh_wire_406[ 8 ];
	assign fresh_wire_193[ 9 ] = fresh_wire_406[ 9 ];
	assign fresh_wire_193[ 10 ] = fresh_wire_406[ 10 ];
	assign fresh_wire_193[ 11 ] = fresh_wire_406[ 11 ];
	assign fresh_wire_193[ 12 ] = fresh_wire_406[ 12 ];
	assign fresh_wire_193[ 13 ] = fresh_wire_406[ 13 ];
	assign fresh_wire_193[ 14 ] = fresh_wire_406[ 14 ];
	assign fresh_wire_193[ 15 ] = fresh_wire_406[ 15 ];
	assign fresh_wire_194[ 0 ] = fresh_wire_1156[ 0 ];
	assign fresh_wire_194[ 1 ] = fresh_wire_1156[ 1 ];
	assign fresh_wire_194[ 2 ] = fresh_wire_1156[ 2 ];
	assign fresh_wire_194[ 3 ] = fresh_wire_1156[ 3 ];
	assign fresh_wire_194[ 4 ] = fresh_wire_1156[ 4 ];
	assign fresh_wire_194[ 5 ] = fresh_wire_1156[ 5 ];
	assign fresh_wire_194[ 6 ] = fresh_wire_1156[ 6 ];
	assign fresh_wire_194[ 7 ] = fresh_wire_1156[ 7 ];
	assign fresh_wire_194[ 8 ] = fresh_wire_1156[ 8 ];
	assign fresh_wire_194[ 9 ] = fresh_wire_1156[ 9 ];
	assign fresh_wire_194[ 10 ] = fresh_wire_1156[ 10 ];
	assign fresh_wire_194[ 11 ] = fresh_wire_1156[ 11 ];
	assign fresh_wire_194[ 12 ] = fresh_wire_1156[ 12 ];
	assign fresh_wire_194[ 13 ] = fresh_wire_1156[ 13 ];
	assign fresh_wire_194[ 14 ] = fresh_wire_1156[ 14 ];
	assign fresh_wire_194[ 15 ] = fresh_wire_1156[ 15 ];
	assign fresh_wire_196[ 0 ] = fresh_wire_406[ 0 ];
	assign fresh_wire_196[ 1 ] = fresh_wire_406[ 1 ];
	assign fresh_wire_196[ 2 ] = fresh_wire_406[ 2 ];
	assign fresh_wire_196[ 3 ] = fresh_wire_406[ 3 ];
	assign fresh_wire_196[ 4 ] = fresh_wire_406[ 4 ];
	assign fresh_wire_196[ 5 ] = fresh_wire_406[ 5 ];
	assign fresh_wire_196[ 6 ] = fresh_wire_406[ 6 ];
	assign fresh_wire_196[ 7 ] = fresh_wire_406[ 7 ];
	assign fresh_wire_196[ 8 ] = fresh_wire_406[ 8 ];
	assign fresh_wire_196[ 9 ] = fresh_wire_406[ 9 ];
	assign fresh_wire_196[ 10 ] = fresh_wire_406[ 10 ];
	assign fresh_wire_196[ 11 ] = fresh_wire_406[ 11 ];
	assign fresh_wire_196[ 12 ] = fresh_wire_406[ 12 ];
	assign fresh_wire_196[ 13 ] = fresh_wire_406[ 13 ];
	assign fresh_wire_196[ 14 ] = fresh_wire_406[ 14 ];
	assign fresh_wire_196[ 15 ] = fresh_wire_406[ 15 ];
	assign fresh_wire_197[ 0 ] = fresh_wire_1157[ 0 ];
	assign fresh_wire_197[ 1 ] = fresh_wire_1157[ 1 ];
	assign fresh_wire_197[ 2 ] = fresh_wire_1157[ 2 ];
	assign fresh_wire_197[ 3 ] = fresh_wire_1157[ 3 ];
	assign fresh_wire_197[ 4 ] = fresh_wire_1157[ 4 ];
	assign fresh_wire_197[ 5 ] = fresh_wire_1157[ 5 ];
	assign fresh_wire_197[ 6 ] = fresh_wire_1157[ 6 ];
	assign fresh_wire_197[ 7 ] = fresh_wire_1157[ 7 ];
	assign fresh_wire_197[ 8 ] = fresh_wire_1157[ 8 ];
	assign fresh_wire_197[ 9 ] = fresh_wire_1157[ 9 ];
	assign fresh_wire_197[ 10 ] = fresh_wire_1157[ 10 ];
	assign fresh_wire_197[ 11 ] = fresh_wire_1157[ 11 ];
	assign fresh_wire_197[ 12 ] = fresh_wire_1157[ 12 ];
	assign fresh_wire_197[ 13 ] = fresh_wire_1157[ 13 ];
	assign fresh_wire_197[ 14 ] = fresh_wire_1157[ 14 ];
	assign fresh_wire_197[ 15 ] = fresh_wire_1157[ 15 ];
	assign fresh_wire_199[ 0 ] = fresh_wire_219[ 0 ];
	assign fresh_wire_200[ 0 ] = fresh_wire_228[ 0 ];
	assign fresh_wire_202[ 0 ] = fresh_wire_376[ 0 ];
	assign fresh_wire_202[ 1 ] = fresh_wire_376[ 1 ];
	assign fresh_wire_203[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_203[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_205[ 0 ] = fresh_wire_373[ 0 ];
	assign fresh_wire_205[ 1 ] = fresh_wire_373[ 1 ];
	assign fresh_wire_206[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_206[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_208[ 0 ] = fresh_wire_666[ 0 ];
	assign fresh_wire_208[ 1 ] = fresh_wire_666[ 1 ];
	assign fresh_wire_209[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_209[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_211[ 0 ] = fresh_wire_166[ 0 ];
	assign fresh_wire_211[ 1 ] = fresh_wire_166[ 1 ];
	assign fresh_wire_211[ 2 ] = fresh_wire_166[ 2 ];
	assign fresh_wire_211[ 3 ] = fresh_wire_166[ 3 ];
	assign fresh_wire_211[ 4 ] = fresh_wire_166[ 4 ];
	assign fresh_wire_211[ 5 ] = fresh_wire_166[ 5 ];
	assign fresh_wire_211[ 6 ] = fresh_wire_166[ 6 ];
	assign fresh_wire_211[ 7 ] = fresh_wire_166[ 7 ];
	assign fresh_wire_211[ 8 ] = fresh_wire_166[ 8 ];
	assign fresh_wire_211[ 9 ] = fresh_wire_166[ 9 ];
	assign fresh_wire_211[ 10 ] = fresh_wire_166[ 10 ];
	assign fresh_wire_211[ 11 ] = fresh_wire_166[ 11 ];
	assign fresh_wire_211[ 12 ] = fresh_wire_166[ 12 ];
	assign fresh_wire_211[ 13 ] = fresh_wire_166[ 13 ];
	assign fresh_wire_211[ 14 ] = fresh_wire_166[ 14 ];
	assign fresh_wire_211[ 15 ] = fresh_wire_166[ 15 ];
	assign fresh_wire_212[ 0 ] = fresh_wire_1158[ 0 ];
	assign fresh_wire_212[ 1 ] = fresh_wire_1158[ 1 ];
	assign fresh_wire_212[ 2 ] = fresh_wire_1158[ 2 ];
	assign fresh_wire_212[ 3 ] = fresh_wire_1158[ 3 ];
	assign fresh_wire_212[ 4 ] = fresh_wire_1158[ 4 ];
	assign fresh_wire_212[ 5 ] = fresh_wire_1158[ 5 ];
	assign fresh_wire_212[ 6 ] = fresh_wire_1158[ 6 ];
	assign fresh_wire_212[ 7 ] = fresh_wire_1158[ 7 ];
	assign fresh_wire_212[ 8 ] = fresh_wire_1158[ 8 ];
	assign fresh_wire_212[ 9 ] = fresh_wire_1158[ 9 ];
	assign fresh_wire_212[ 10 ] = fresh_wire_1158[ 10 ];
	assign fresh_wire_212[ 11 ] = fresh_wire_1158[ 11 ];
	assign fresh_wire_212[ 12 ] = fresh_wire_1158[ 12 ];
	assign fresh_wire_212[ 13 ] = fresh_wire_1158[ 13 ];
	assign fresh_wire_212[ 14 ] = fresh_wire_1158[ 14 ];
	assign fresh_wire_212[ 15 ] = fresh_wire_1158[ 15 ];
	assign fresh_wire_214[ 0 ] = fresh_wire_422[ 0 ];
	assign fresh_wire_215[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_217[ 0 ] = fresh_wire_430[ 0 ];
	assign fresh_wire_218[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_220[ 0 ] = fresh_wire_678[ 0 ];
	assign fresh_wire_221[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_223[ 0 ] = fresh_wire_286[ 0 ];
	assign fresh_wire_224[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_226[ 0 ] = fresh_wire_402[ 0 ];
	assign fresh_wire_226[ 1 ] = fresh_wire_402[ 1 ];
	assign fresh_wire_227[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_227[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_229[ 0 ] = fresh_wire_430[ 0 ];
	assign fresh_wire_230[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_232[ 0 ] = fresh_wire_426[ 0 ];
	assign fresh_wire_233[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_235[ 0 ] = fresh_wire_402[ 0 ];
	assign fresh_wire_235[ 1 ] = fresh_wire_402[ 1 ];
	assign fresh_wire_236[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_236[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_238[ 0 ] = fresh_wire_363[ 0 ];
	assign fresh_wire_239[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_241[ 0 ] = fresh_wire_398[ 0 ];
	assign fresh_wire_242[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_244[ 0 ] = fresh_wire_402[ 0 ];
	assign fresh_wire_244[ 1 ] = fresh_wire_402[ 1 ];
	assign fresh_wire_245[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_245[ 1 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_247[ 0 ] = fresh_wire_373[ 0 ];
	assign fresh_wire_247[ 1 ] = fresh_wire_373[ 1 ];
	assign fresh_wire_248[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_248[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_250[ 0 ] = fresh_wire_198[ 0 ];
	assign fresh_wire_250[ 1 ] = fresh_wire_198[ 1 ];
	assign fresh_wire_250[ 2 ] = fresh_wire_198[ 2 ];
	assign fresh_wire_250[ 3 ] = fresh_wire_198[ 3 ];
	assign fresh_wire_250[ 4 ] = fresh_wire_198[ 4 ];
	assign fresh_wire_250[ 5 ] = fresh_wire_198[ 5 ];
	assign fresh_wire_250[ 6 ] = fresh_wire_198[ 6 ];
	assign fresh_wire_250[ 7 ] = fresh_wire_198[ 7 ];
	assign fresh_wire_250[ 8 ] = fresh_wire_198[ 8 ];
	assign fresh_wire_250[ 9 ] = fresh_wire_198[ 9 ];
	assign fresh_wire_250[ 10 ] = fresh_wire_198[ 10 ];
	assign fresh_wire_250[ 11 ] = fresh_wire_198[ 11 ];
	assign fresh_wire_250[ 12 ] = fresh_wire_198[ 12 ];
	assign fresh_wire_250[ 13 ] = fresh_wire_198[ 13 ];
	assign fresh_wire_250[ 14 ] = fresh_wire_198[ 14 ];
	assign fresh_wire_250[ 15 ] = fresh_wire_198[ 15 ];
	assign fresh_wire_251[ 0 ] = fresh_wire_1159[ 0 ];
	assign fresh_wire_251[ 1 ] = fresh_wire_1159[ 1 ];
	assign fresh_wire_251[ 2 ] = fresh_wire_1159[ 2 ];
	assign fresh_wire_251[ 3 ] = fresh_wire_1159[ 3 ];
	assign fresh_wire_251[ 4 ] = fresh_wire_1159[ 4 ];
	assign fresh_wire_251[ 5 ] = fresh_wire_1159[ 5 ];
	assign fresh_wire_251[ 6 ] = fresh_wire_1159[ 6 ];
	assign fresh_wire_251[ 7 ] = fresh_wire_1159[ 7 ];
	assign fresh_wire_251[ 8 ] = fresh_wire_1159[ 8 ];
	assign fresh_wire_251[ 9 ] = fresh_wire_1159[ 9 ];
	assign fresh_wire_251[ 10 ] = fresh_wire_1159[ 10 ];
	assign fresh_wire_251[ 11 ] = fresh_wire_1159[ 11 ];
	assign fresh_wire_251[ 12 ] = fresh_wire_1159[ 12 ];
	assign fresh_wire_251[ 13 ] = fresh_wire_1159[ 13 ];
	assign fresh_wire_251[ 14 ] = fresh_wire_1159[ 14 ];
	assign fresh_wire_251[ 15 ] = fresh_wire_1159[ 15 ];
	assign fresh_wire_253[ 0 ] = fresh_wire_894[ 0 ];
	assign fresh_wire_254[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_256[ 0 ] = fresh_wire_394[ 0 ];
	assign fresh_wire_257[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_259[ 0 ] = fresh_wire_414[ 0 ];
	assign fresh_wire_259[ 1 ] = fresh_wire_414[ 1 ];
	assign fresh_wire_259[ 2 ] = fresh_wire_414[ 2 ];
	assign fresh_wire_259[ 3 ] = fresh_wire_414[ 3 ];
	assign fresh_wire_259[ 4 ] = fresh_wire_414[ 4 ];
	assign fresh_wire_259[ 5 ] = fresh_wire_414[ 5 ];
	assign fresh_wire_259[ 6 ] = fresh_wire_414[ 6 ];
	assign fresh_wire_259[ 7 ] = fresh_wire_414[ 7 ];
	assign fresh_wire_259[ 8 ] = fresh_wire_414[ 8 ];
	assign fresh_wire_259[ 9 ] = fresh_wire_414[ 9 ];
	assign fresh_wire_259[ 10 ] = fresh_wire_414[ 10 ];
	assign fresh_wire_259[ 11 ] = fresh_wire_414[ 11 ];
	assign fresh_wire_259[ 12 ] = fresh_wire_414[ 12 ];
	assign fresh_wire_259[ 13 ] = fresh_wire_414[ 13 ];
	assign fresh_wire_259[ 14 ] = fresh_wire_414[ 14 ];
	assign fresh_wire_259[ 15 ] = fresh_wire_414[ 15 ];
	assign fresh_wire_260[ 0 ] = fresh_wire_1161[ 0 ];
	assign fresh_wire_260[ 1 ] = fresh_wire_1161[ 1 ];
	assign fresh_wire_260[ 2 ] = fresh_wire_1161[ 2 ];
	assign fresh_wire_260[ 3 ] = fresh_wire_1161[ 3 ];
	assign fresh_wire_260[ 4 ] = fresh_wire_1161[ 4 ];
	assign fresh_wire_260[ 5 ] = fresh_wire_1161[ 5 ];
	assign fresh_wire_260[ 6 ] = fresh_wire_1161[ 6 ];
	assign fresh_wire_260[ 7 ] = fresh_wire_1161[ 7 ];
	assign fresh_wire_260[ 8 ] = fresh_wire_1161[ 8 ];
	assign fresh_wire_260[ 9 ] = fresh_wire_1161[ 9 ];
	assign fresh_wire_260[ 10 ] = fresh_wire_1161[ 10 ];
	assign fresh_wire_260[ 11 ] = fresh_wire_1161[ 11 ];
	assign fresh_wire_260[ 12 ] = fresh_wire_1161[ 12 ];
	assign fresh_wire_260[ 13 ] = fresh_wire_1161[ 13 ];
	assign fresh_wire_260[ 14 ] = fresh_wire_1161[ 14 ];
	assign fresh_wire_260[ 15 ] = fresh_wire_1161[ 15 ];
	assign fresh_wire_262[ 0 ] = fresh_wire_410[ 0 ];
	assign fresh_wire_262[ 1 ] = fresh_wire_410[ 1 ];
	assign fresh_wire_262[ 2 ] = fresh_wire_410[ 2 ];
	assign fresh_wire_262[ 3 ] = fresh_wire_410[ 3 ];
	assign fresh_wire_262[ 4 ] = fresh_wire_410[ 4 ];
	assign fresh_wire_262[ 5 ] = fresh_wire_410[ 5 ];
	assign fresh_wire_262[ 6 ] = fresh_wire_410[ 6 ];
	assign fresh_wire_262[ 7 ] = fresh_wire_410[ 7 ];
	assign fresh_wire_262[ 8 ] = fresh_wire_410[ 8 ];
	assign fresh_wire_262[ 9 ] = fresh_wire_410[ 9 ];
	assign fresh_wire_262[ 10 ] = fresh_wire_410[ 10 ];
	assign fresh_wire_262[ 11 ] = fresh_wire_410[ 11 ];
	assign fresh_wire_262[ 12 ] = fresh_wire_410[ 12 ];
	assign fresh_wire_262[ 13 ] = fresh_wire_410[ 13 ];
	assign fresh_wire_262[ 14 ] = fresh_wire_410[ 14 ];
	assign fresh_wire_262[ 15 ] = fresh_wire_410[ 15 ];
	assign fresh_wire_263[ 0 ] = fresh_wire_1161[ 0 ];
	assign fresh_wire_263[ 1 ] = fresh_wire_1161[ 1 ];
	assign fresh_wire_263[ 2 ] = fresh_wire_1161[ 2 ];
	assign fresh_wire_263[ 3 ] = fresh_wire_1161[ 3 ];
	assign fresh_wire_263[ 4 ] = fresh_wire_1161[ 4 ];
	assign fresh_wire_263[ 5 ] = fresh_wire_1161[ 5 ];
	assign fresh_wire_263[ 6 ] = fresh_wire_1161[ 6 ];
	assign fresh_wire_263[ 7 ] = fresh_wire_1161[ 7 ];
	assign fresh_wire_263[ 8 ] = fresh_wire_1161[ 8 ];
	assign fresh_wire_263[ 9 ] = fresh_wire_1161[ 9 ];
	assign fresh_wire_263[ 10 ] = fresh_wire_1161[ 10 ];
	assign fresh_wire_263[ 11 ] = fresh_wire_1161[ 11 ];
	assign fresh_wire_263[ 12 ] = fresh_wire_1161[ 12 ];
	assign fresh_wire_263[ 13 ] = fresh_wire_1161[ 13 ];
	assign fresh_wire_263[ 14 ] = fresh_wire_1161[ 14 ];
	assign fresh_wire_263[ 15 ] = fresh_wire_1161[ 15 ];
	assign fresh_wire_265[ 0 ] = fresh_wire_195[ 0 ];
	assign fresh_wire_265[ 1 ] = fresh_wire_195[ 1 ];
	assign fresh_wire_265[ 2 ] = fresh_wire_195[ 2 ];
	assign fresh_wire_265[ 3 ] = fresh_wire_195[ 3 ];
	assign fresh_wire_265[ 4 ] = fresh_wire_195[ 4 ];
	assign fresh_wire_265[ 5 ] = fresh_wire_195[ 5 ];
	assign fresh_wire_265[ 6 ] = fresh_wire_195[ 6 ];
	assign fresh_wire_265[ 7 ] = fresh_wire_195[ 7 ];
	assign fresh_wire_265[ 8 ] = fresh_wire_195[ 8 ];
	assign fresh_wire_265[ 9 ] = fresh_wire_195[ 9 ];
	assign fresh_wire_265[ 10 ] = fresh_wire_195[ 10 ];
	assign fresh_wire_265[ 11 ] = fresh_wire_195[ 11 ];
	assign fresh_wire_265[ 12 ] = fresh_wire_195[ 12 ];
	assign fresh_wire_265[ 13 ] = fresh_wire_195[ 13 ];
	assign fresh_wire_265[ 14 ] = fresh_wire_195[ 14 ];
	assign fresh_wire_265[ 15 ] = fresh_wire_195[ 15 ];
	assign fresh_wire_266[ 0 ] = fresh_wire_1160[ 0 ];
	assign fresh_wire_266[ 1 ] = fresh_wire_1160[ 1 ];
	assign fresh_wire_266[ 2 ] = fresh_wire_1160[ 2 ];
	assign fresh_wire_266[ 3 ] = fresh_wire_1160[ 3 ];
	assign fresh_wire_266[ 4 ] = fresh_wire_1160[ 4 ];
	assign fresh_wire_266[ 5 ] = fresh_wire_1160[ 5 ];
	assign fresh_wire_266[ 6 ] = fresh_wire_1160[ 6 ];
	assign fresh_wire_266[ 7 ] = fresh_wire_1160[ 7 ];
	assign fresh_wire_266[ 8 ] = fresh_wire_1160[ 8 ];
	assign fresh_wire_266[ 9 ] = fresh_wire_1160[ 9 ];
	assign fresh_wire_266[ 10 ] = fresh_wire_1160[ 10 ];
	assign fresh_wire_266[ 11 ] = fresh_wire_1160[ 11 ];
	assign fresh_wire_266[ 12 ] = fresh_wire_1160[ 12 ];
	assign fresh_wire_266[ 13 ] = fresh_wire_1160[ 13 ];
	assign fresh_wire_266[ 14 ] = fresh_wire_1160[ 14 ];
	assign fresh_wire_266[ 15 ] = fresh_wire_1160[ 15 ];
	assign fresh_wire_268[ 0 ] = fresh_wire_204[ 0 ];
	assign fresh_wire_270[ 0 ] = fresh_wire_269[ 0 ];
	assign fresh_wire_271[ 0 ] = fresh_wire_274[ 0 ];
	assign fresh_wire_273[ 0 ] = fresh_wire_207[ 0 ];
	assign fresh_wire_275[ 0 ] = fresh_wire_272[ 0 ];
	assign fresh_wire_277[ 0 ] = fresh_wire_276[ 0 ];
	assign fresh_wire_278[ 0 ] = fresh_wire_281[ 0 ];
	assign fresh_wire_280[ 0 ] = fresh_wire_210[ 0 ];
	assign fresh_wire_282[ 0 ] = fresh_wire_279[ 0 ];
	assign fresh_wire_284[ 0 ] = fresh_wire_283[ 0 ];
	assign fresh_wire_285[ 0 ] = fresh_wire_288[ 0 ];
	assign fresh_wire_287[ 0 ] = fresh_wire_213[ 0 ];
	assign fresh_wire_289[ 0 ] = fresh_wire_237[ 0 ];
	assign fresh_wire_291[ 0 ] = fresh_wire_290[ 0 ];
	assign fresh_wire_292[ 0 ] = fresh_wire_1175[ 0 ];
	assign fresh_wire_294[ 0 ] = fresh_wire_293[ 0 ];
	assign fresh_wire_296[ 0 ] = fresh_wire_295[ 0 ];
	assign fresh_wire_297[ 0 ] = fresh_wire_300[ 0 ];
	assign fresh_wire_299[ 0 ] = fresh_wire_240[ 0 ];
	assign fresh_wire_301[ 0 ] = fresh_wire_228[ 0 ];
	assign fresh_wire_303[ 0 ] = fresh_wire_302[ 0 ];
	assign fresh_wire_304[ 0 ] = fresh_wire_1176[ 0 ];
	assign fresh_wire_306[ 0 ] = fresh_wire_305[ 0 ];
	assign fresh_wire_308[ 0 ] = fresh_wire_307[ 0 ];
	assign fresh_wire_309[ 0 ] = fresh_wire_312[ 0 ];
	assign fresh_wire_311[ 0 ] = fresh_wire_366[ 0 ];
	assign fresh_wire_313[ 0 ] = fresh_wire_228[ 0 ];
	assign fresh_wire_315[ 0 ] = fresh_wire_314[ 0 ];
	assign fresh_wire_316[ 0 ] = fresh_wire_319[ 0 ];
	assign fresh_wire_318[ 0 ] = fresh_wire_267[ 0 ];
	assign fresh_wire_320[ 0 ] = fresh_wire_1177[ 0 ];
	assign fresh_wire_321[ 0 ] = fresh_wire_324[ 0 ];
	assign fresh_wire_323[ 0 ] = fresh_wire_240[ 0 ];
	assign fresh_wire_325[ 0 ] = fresh_wire_246[ 0 ];
	assign fresh_wire_327[ 0 ] = fresh_wire_326[ 0 ];
	assign fresh_wire_328[ 0 ] = fresh_wire_1178[ 0 ];
	assign fresh_wire_330[ 0 ] = fresh_wire_204[ 0 ];
	assign fresh_wire_332[ 0 ] = fresh_wire_331[ 0 ];
	assign fresh_wire_333[ 0 ] = fresh_wire_336[ 0 ];
	assign fresh_wire_335[ 0 ] = fresh_wire_207[ 0 ];
	assign fresh_wire_337[ 0 ] = fresh_wire_334[ 0 ];
	assign fresh_wire_339[ 0 ] = fresh_wire_338[ 0 ];
	assign fresh_wire_340[ 0 ] = fresh_wire_343[ 0 ];
	assign fresh_wire_342[ 0 ] = fresh_wire_210[ 0 ];
	assign fresh_wire_344[ 0 ] = fresh_wire_341[ 0 ];
	assign fresh_wire_346[ 0 ] = fresh_wire_345[ 0 ];
	assign fresh_wire_347[ 0 ] = fresh_wire_350[ 0 ];
	assign fresh_wire_349[ 0 ] = fresh_wire_252[ 0 ];
	assign fresh_wire_351[ 0 ] = fresh_wire_255[ 0 ];
	assign fresh_wire_353[ 0 ] = fresh_wire_352[ 0 ];
	assign fresh_wire_354[ 0 ] = fresh_wire_1179[ 0 ];
	assign fresh_wire_356[ 0 ] = fresh_wire_363[ 0 ];
	assign fresh_wire_358[ 0 ] = fresh_wire_1180[ 0 ];
	assign fresh_wire_359[ 0 ] = fresh_wire_357[ 0 ];
	assign fresh_wire_361[ 0 ] = fresh_wire_171[ 0 ];
	assign fresh_wire_361[ 1 ] = fresh_wire_171[ 1 ];
	assign fresh_wire_361[ 2 ] = fresh_wire_171[ 2 ];
	assign fresh_wire_361[ 3 ] = fresh_wire_171[ 3 ];
	assign fresh_wire_361[ 4 ] = fresh_wire_171[ 4 ];
	assign fresh_wire_361[ 5 ] = fresh_wire_171[ 5 ];
	assign fresh_wire_361[ 6 ] = fresh_wire_171[ 6 ];
	assign fresh_wire_361[ 7 ] = fresh_wire_171[ 7 ];
	assign fresh_wire_361[ 8 ] = fresh_wire_171[ 8 ];
	assign fresh_wire_361[ 9 ] = fresh_wire_171[ 9 ];
	assign fresh_wire_361[ 10 ] = fresh_wire_171[ 10 ];
	assign fresh_wire_361[ 11 ] = fresh_wire_171[ 11 ];
	assign fresh_wire_361[ 12 ] = fresh_wire_171[ 12 ];
	assign fresh_wire_361[ 13 ] = fresh_wire_171[ 13 ];
	assign fresh_wire_361[ 14 ] = fresh_wire_171[ 14 ];
	assign fresh_wire_361[ 15 ] = fresh_wire_171[ 15 ];
	assign fresh_wire_362[ 0 ] = fresh_wire_1162[ 0 ];
	assign fresh_wire_362[ 1 ] = fresh_wire_1162[ 1 ];
	assign fresh_wire_362[ 2 ] = fresh_wire_1162[ 2 ];
	assign fresh_wire_362[ 3 ] = fresh_wire_1162[ 3 ];
	assign fresh_wire_362[ 4 ] = fresh_wire_1162[ 4 ];
	assign fresh_wire_362[ 5 ] = fresh_wire_1162[ 5 ];
	assign fresh_wire_362[ 6 ] = fresh_wire_1162[ 6 ];
	assign fresh_wire_362[ 7 ] = fresh_wire_1162[ 7 ];
	assign fresh_wire_362[ 8 ] = fresh_wire_1162[ 8 ];
	assign fresh_wire_362[ 9 ] = fresh_wire_1162[ 9 ];
	assign fresh_wire_362[ 10 ] = fresh_wire_1162[ 10 ];
	assign fresh_wire_362[ 11 ] = fresh_wire_1162[ 11 ];
	assign fresh_wire_362[ 12 ] = fresh_wire_1162[ 12 ];
	assign fresh_wire_362[ 13 ] = fresh_wire_1162[ 13 ];
	assign fresh_wire_362[ 14 ] = fresh_wire_1162[ 14 ];
	assign fresh_wire_362[ 15 ] = fresh_wire_1162[ 15 ];
	assign fresh_wire_364[ 0 ] = fresh_wire_189[ 0 ];
	assign fresh_wire_364[ 1 ] = fresh_wire_189[ 1 ];
	assign fresh_wire_364[ 2 ] = fresh_wire_189[ 2 ];
	assign fresh_wire_364[ 3 ] = fresh_wire_189[ 3 ];
	assign fresh_wire_364[ 4 ] = fresh_wire_189[ 4 ];
	assign fresh_wire_364[ 5 ] = fresh_wire_189[ 5 ];
	assign fresh_wire_364[ 6 ] = fresh_wire_189[ 6 ];
	assign fresh_wire_364[ 7 ] = fresh_wire_189[ 7 ];
	assign fresh_wire_364[ 8 ] = fresh_wire_189[ 8 ];
	assign fresh_wire_364[ 9 ] = fresh_wire_189[ 9 ];
	assign fresh_wire_364[ 10 ] = fresh_wire_189[ 10 ];
	assign fresh_wire_364[ 11 ] = fresh_wire_189[ 11 ];
	assign fresh_wire_364[ 12 ] = fresh_wire_189[ 12 ];
	assign fresh_wire_364[ 13 ] = fresh_wire_189[ 13 ];
	assign fresh_wire_364[ 14 ] = fresh_wire_189[ 14 ];
	assign fresh_wire_364[ 15 ] = fresh_wire_189[ 15 ];
	assign fresh_wire_365[ 0 ] = fresh_wire_1160[ 0 ];
	assign fresh_wire_365[ 1 ] = fresh_wire_1160[ 1 ];
	assign fresh_wire_365[ 2 ] = fresh_wire_1160[ 2 ];
	assign fresh_wire_365[ 3 ] = fresh_wire_1160[ 3 ];
	assign fresh_wire_365[ 4 ] = fresh_wire_1160[ 4 ];
	assign fresh_wire_365[ 5 ] = fresh_wire_1160[ 5 ];
	assign fresh_wire_365[ 6 ] = fresh_wire_1160[ 6 ];
	assign fresh_wire_365[ 7 ] = fresh_wire_1160[ 7 ];
	assign fresh_wire_365[ 8 ] = fresh_wire_1160[ 8 ];
	assign fresh_wire_365[ 9 ] = fresh_wire_1160[ 9 ];
	assign fresh_wire_365[ 10 ] = fresh_wire_1160[ 10 ];
	assign fresh_wire_365[ 11 ] = fresh_wire_1160[ 11 ];
	assign fresh_wire_365[ 12 ] = fresh_wire_1160[ 12 ];
	assign fresh_wire_365[ 13 ] = fresh_wire_1160[ 13 ];
	assign fresh_wire_365[ 14 ] = fresh_wire_1160[ 14 ];
	assign fresh_wire_365[ 15 ] = fresh_wire_1160[ 15 ];
	assign fresh_wire_367[ 0 ] = fresh_wire_430[ 0 ];
	assign fresh_wire_369[ 0 ] = fresh_wire_360[ 0 ];
	assign fresh_wire_371[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_372[ 0 ] = fresh_wire_402[ 0 ];
	assign fresh_wire_372[ 1 ] = fresh_wire_402[ 1 ];
	assign fresh_wire_374[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_375[ 0 ] = fresh_wire_373[ 0 ];
	assign fresh_wire_375[ 1 ] = fresh_wire_373[ 1 ];
	assign fresh_wire_377[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_378[ 0 ] = fresh_wire_878[ 0 ];
	assign fresh_wire_378[ 1 ] = fresh_wire_878[ 1 ];
	assign fresh_wire_378[ 2 ] = fresh_wire_878[ 2 ];
	assign fresh_wire_378[ 3 ] = fresh_wire_878[ 3 ];
	assign fresh_wire_378[ 4 ] = fresh_wire_878[ 4 ];
	assign fresh_wire_378[ 5 ] = fresh_wire_878[ 5 ];
	assign fresh_wire_378[ 6 ] = fresh_wire_878[ 6 ];
	assign fresh_wire_378[ 7 ] = fresh_wire_878[ 7 ];
	assign fresh_wire_378[ 8 ] = fresh_wire_878[ 8 ];
	assign fresh_wire_378[ 9 ] = fresh_wire_878[ 9 ];
	assign fresh_wire_378[ 10 ] = fresh_wire_878[ 10 ];
	assign fresh_wire_378[ 11 ] = fresh_wire_878[ 11 ];
	assign fresh_wire_378[ 12 ] = fresh_wire_878[ 12 ];
	assign fresh_wire_378[ 13 ] = fresh_wire_878[ 13 ];
	assign fresh_wire_378[ 14 ] = fresh_wire_878[ 14 ];
	assign fresh_wire_378[ 15 ] = fresh_wire_878[ 15 ];
	assign fresh_wire_380[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_381[ 0 ] = fresh_wire_455[ 0 ];
	assign fresh_wire_383[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_384[ 0 ] = fresh_wire_1153[ 0 ];
	assign fresh_wire_385[ 0 ] = fresh_wire_451[ 0 ];
	assign fresh_wire_387[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_388[ 0 ] = fresh_wire_1153[ 0 ];
	assign fresh_wire_389[ 0 ] = fresh_wire_443[ 0 ];
	assign fresh_wire_391[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_392[ 0 ] = fresh_wire_1153[ 0 ];
	assign fresh_wire_393[ 0 ] = fresh_wire_535[ 0 ];
	assign fresh_wire_395[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_396[ 0 ] = fresh_wire_1153[ 0 ];
	assign fresh_wire_397[ 0 ] = fresh_wire_511[ 0 ];
	assign fresh_wire_399[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_400[ 0 ] = fresh_wire_1153[ 0 ];
	assign fresh_wire_401[ 0 ] = fresh_wire_495[ 0 ];
	assign fresh_wire_401[ 1 ] = fresh_wire_495[ 1 ];
	assign fresh_wire_403[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_404[ 0 ] = fresh_wire_1153[ 0 ];
	assign fresh_wire_405[ 0 ] = fresh_wire_471[ 0 ];
	assign fresh_wire_405[ 1 ] = fresh_wire_471[ 1 ];
	assign fresh_wire_405[ 2 ] = fresh_wire_471[ 2 ];
	assign fresh_wire_405[ 3 ] = fresh_wire_471[ 3 ];
	assign fresh_wire_405[ 4 ] = fresh_wire_471[ 4 ];
	assign fresh_wire_405[ 5 ] = fresh_wire_471[ 5 ];
	assign fresh_wire_405[ 6 ] = fresh_wire_471[ 6 ];
	assign fresh_wire_405[ 7 ] = fresh_wire_471[ 7 ];
	assign fresh_wire_405[ 8 ] = fresh_wire_471[ 8 ];
	assign fresh_wire_405[ 9 ] = fresh_wire_471[ 9 ];
	assign fresh_wire_405[ 10 ] = fresh_wire_471[ 10 ];
	assign fresh_wire_405[ 11 ] = fresh_wire_471[ 11 ];
	assign fresh_wire_405[ 12 ] = fresh_wire_471[ 12 ];
	assign fresh_wire_405[ 13 ] = fresh_wire_471[ 13 ];
	assign fresh_wire_405[ 14 ] = fresh_wire_471[ 14 ];
	assign fresh_wire_405[ 15 ] = fresh_wire_471[ 15 ];
	assign fresh_wire_407[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_408[ 0 ] = fresh_wire_1153[ 0 ];
	assign fresh_wire_409[ 0 ] = fresh_wire_571[ 0 ];
	assign fresh_wire_409[ 1 ] = fresh_wire_571[ 1 ];
	assign fresh_wire_409[ 2 ] = fresh_wire_571[ 2 ];
	assign fresh_wire_409[ 3 ] = fresh_wire_571[ 3 ];
	assign fresh_wire_409[ 4 ] = fresh_wire_571[ 4 ];
	assign fresh_wire_409[ 5 ] = fresh_wire_571[ 5 ];
	assign fresh_wire_409[ 6 ] = fresh_wire_571[ 6 ];
	assign fresh_wire_409[ 7 ] = fresh_wire_571[ 7 ];
	assign fresh_wire_409[ 8 ] = fresh_wire_571[ 8 ];
	assign fresh_wire_409[ 9 ] = fresh_wire_571[ 9 ];
	assign fresh_wire_409[ 10 ] = fresh_wire_571[ 10 ];
	assign fresh_wire_409[ 11 ] = fresh_wire_571[ 11 ];
	assign fresh_wire_409[ 12 ] = fresh_wire_571[ 12 ];
	assign fresh_wire_409[ 13 ] = fresh_wire_571[ 13 ];
	assign fresh_wire_409[ 14 ] = fresh_wire_571[ 14 ];
	assign fresh_wire_409[ 15 ] = fresh_wire_571[ 15 ];
	assign fresh_wire_411[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_412[ 0 ] = fresh_wire_1153[ 0 ];
	assign fresh_wire_413[ 0 ] = fresh_wire_559[ 0 ];
	assign fresh_wire_413[ 1 ] = fresh_wire_559[ 1 ];
	assign fresh_wire_413[ 2 ] = fresh_wire_559[ 2 ];
	assign fresh_wire_413[ 3 ] = fresh_wire_559[ 3 ];
	assign fresh_wire_413[ 4 ] = fresh_wire_559[ 4 ];
	assign fresh_wire_413[ 5 ] = fresh_wire_559[ 5 ];
	assign fresh_wire_413[ 6 ] = fresh_wire_559[ 6 ];
	assign fresh_wire_413[ 7 ] = fresh_wire_559[ 7 ];
	assign fresh_wire_413[ 8 ] = fresh_wire_559[ 8 ];
	assign fresh_wire_413[ 9 ] = fresh_wire_559[ 9 ];
	assign fresh_wire_413[ 10 ] = fresh_wire_559[ 10 ];
	assign fresh_wire_413[ 11 ] = fresh_wire_559[ 11 ];
	assign fresh_wire_413[ 12 ] = fresh_wire_559[ 12 ];
	assign fresh_wire_413[ 13 ] = fresh_wire_559[ 13 ];
	assign fresh_wire_413[ 14 ] = fresh_wire_559[ 14 ];
	assign fresh_wire_413[ 15 ] = fresh_wire_559[ 15 ];
	assign fresh_wire_415[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_416[ 0 ] = fresh_wire_1153[ 0 ];
	assign fresh_wire_417[ 0 ] = fresh_wire_547[ 0 ];
	assign fresh_wire_417[ 1 ] = fresh_wire_547[ 1 ];
	assign fresh_wire_417[ 2 ] = fresh_wire_547[ 2 ];
	assign fresh_wire_417[ 3 ] = fresh_wire_547[ 3 ];
	assign fresh_wire_417[ 4 ] = fresh_wire_547[ 4 ];
	assign fresh_wire_417[ 5 ] = fresh_wire_547[ 5 ];
	assign fresh_wire_417[ 6 ] = fresh_wire_547[ 6 ];
	assign fresh_wire_417[ 7 ] = fresh_wire_547[ 7 ];
	assign fresh_wire_417[ 8 ] = fresh_wire_547[ 8 ];
	assign fresh_wire_417[ 9 ] = fresh_wire_547[ 9 ];
	assign fresh_wire_417[ 10 ] = fresh_wire_547[ 10 ];
	assign fresh_wire_417[ 11 ] = fresh_wire_547[ 11 ];
	assign fresh_wire_417[ 12 ] = fresh_wire_547[ 12 ];
	assign fresh_wire_417[ 13 ] = fresh_wire_547[ 13 ];
	assign fresh_wire_417[ 14 ] = fresh_wire_547[ 14 ];
	assign fresh_wire_417[ 15 ] = fresh_wire_547[ 15 ];
	assign fresh_wire_419[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_420[ 0 ] = fresh_wire_1153[ 0 ];
	assign fresh_wire_421[ 0 ] = fresh_wire_591[ 0 ];
	assign fresh_wire_423[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_424[ 0 ] = fresh_wire_1153[ 0 ];
	assign fresh_wire_425[ 0 ] = fresh_wire_579[ 0 ];
	assign fresh_wire_427[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_428[ 0 ] = fresh_wire_1153[ 0 ];
	assign fresh_wire_429[ 0 ] = fresh_wire_368[ 0 ];
	assign fresh_wire_431[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_432[ 0 ] = fresh_wire_1153[ 0 ];
	assign fresh_wire_433[ 0 ] = fresh_wire_414[ 0 ];
	assign fresh_wire_433[ 1 ] = fresh_wire_414[ 1 ];
	assign fresh_wire_433[ 2 ] = fresh_wire_414[ 2 ];
	assign fresh_wire_433[ 3 ] = fresh_wire_414[ 3 ];
	assign fresh_wire_433[ 4 ] = fresh_wire_414[ 4 ];
	assign fresh_wire_433[ 5 ] = fresh_wire_414[ 5 ];
	assign fresh_wire_433[ 6 ] = fresh_wire_414[ 6 ];
	assign fresh_wire_433[ 7 ] = fresh_wire_414[ 7 ];
	assign fresh_wire_433[ 8 ] = fresh_wire_414[ 8 ];
	assign fresh_wire_433[ 9 ] = fresh_wire_414[ 9 ];
	assign fresh_wire_433[ 10 ] = fresh_wire_414[ 10 ];
	assign fresh_wire_433[ 11 ] = fresh_wire_414[ 11 ];
	assign fresh_wire_433[ 12 ] = fresh_wire_414[ 12 ];
	assign fresh_wire_433[ 13 ] = fresh_wire_414[ 13 ];
	assign fresh_wire_433[ 14 ] = fresh_wire_414[ 14 ];
	assign fresh_wire_433[ 15 ] = fresh_wire_414[ 15 ];
	assign fresh_wire_434[ 0 ] = fresh_wire_410[ 0 ];
	assign fresh_wire_434[ 1 ] = fresh_wire_410[ 1 ];
	assign fresh_wire_434[ 2 ] = fresh_wire_410[ 2 ];
	assign fresh_wire_434[ 3 ] = fresh_wire_410[ 3 ];
	assign fresh_wire_434[ 4 ] = fresh_wire_410[ 4 ];
	assign fresh_wire_434[ 5 ] = fresh_wire_410[ 5 ];
	assign fresh_wire_434[ 6 ] = fresh_wire_410[ 6 ];
	assign fresh_wire_434[ 7 ] = fresh_wire_410[ 7 ];
	assign fresh_wire_434[ 8 ] = fresh_wire_410[ 8 ];
	assign fresh_wire_434[ 9 ] = fresh_wire_410[ 9 ];
	assign fresh_wire_434[ 10 ] = fresh_wire_410[ 10 ];
	assign fresh_wire_434[ 11 ] = fresh_wire_410[ 11 ];
	assign fresh_wire_434[ 12 ] = fresh_wire_410[ 12 ];
	assign fresh_wire_434[ 13 ] = fresh_wire_410[ 13 ];
	assign fresh_wire_434[ 14 ] = fresh_wire_410[ 14 ];
	assign fresh_wire_434[ 15 ] = fresh_wire_410[ 15 ];
	assign fresh_wire_436[ 0 ] = fresh_wire_219[ 0 ];
	assign fresh_wire_437[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_438[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_440[ 0 ] = fresh_wire_249[ 0 ];
	assign fresh_wire_441[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_442[ 0 ] = fresh_wire_439[ 0 ];
	assign fresh_wire_444[ 0 ] = fresh_wire_219[ 0 ];
	assign fresh_wire_445[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_446[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_448[ 0 ] = fresh_wire_348[ 0 ];
	assign fresh_wire_449[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_450[ 0 ] = fresh_wire_447[ 0 ];
	assign fresh_wire_452[ 0 ] = fresh_wire_219[ 0 ];
	assign fresh_wire_453[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_454[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_456[ 0 ] = fresh_wire_355[ 0 ];
	assign fresh_wire_457[ 0 ] = fresh_wire_406[ 0 ];
	assign fresh_wire_457[ 1 ] = fresh_wire_406[ 1 ];
	assign fresh_wire_457[ 2 ] = fresh_wire_406[ 2 ];
	assign fresh_wire_457[ 3 ] = fresh_wire_406[ 3 ];
	assign fresh_wire_457[ 4 ] = fresh_wire_406[ 4 ];
	assign fresh_wire_457[ 5 ] = fresh_wire_406[ 5 ];
	assign fresh_wire_457[ 6 ] = fresh_wire_406[ 6 ];
	assign fresh_wire_457[ 7 ] = fresh_wire_406[ 7 ];
	assign fresh_wire_457[ 8 ] = fresh_wire_406[ 8 ];
	assign fresh_wire_457[ 9 ] = fresh_wire_406[ 9 ];
	assign fresh_wire_457[ 10 ] = fresh_wire_406[ 10 ];
	assign fresh_wire_457[ 11 ] = fresh_wire_406[ 11 ];
	assign fresh_wire_457[ 12 ] = fresh_wire_406[ 12 ];
	assign fresh_wire_457[ 13 ] = fresh_wire_406[ 13 ];
	assign fresh_wire_457[ 14 ] = fresh_wire_406[ 14 ];
	assign fresh_wire_457[ 15 ] = fresh_wire_406[ 15 ];
	assign fresh_wire_458[ 0 ] = fresh_wire_192[ 0 ];
	assign fresh_wire_458[ 1 ] = fresh_wire_192[ 1 ];
	assign fresh_wire_458[ 2 ] = fresh_wire_192[ 2 ];
	assign fresh_wire_458[ 3 ] = fresh_wire_192[ 3 ];
	assign fresh_wire_458[ 4 ] = fresh_wire_192[ 4 ];
	assign fresh_wire_458[ 5 ] = fresh_wire_192[ 5 ];
	assign fresh_wire_458[ 6 ] = fresh_wire_192[ 6 ];
	assign fresh_wire_458[ 7 ] = fresh_wire_192[ 7 ];
	assign fresh_wire_458[ 8 ] = fresh_wire_192[ 8 ];
	assign fresh_wire_458[ 9 ] = fresh_wire_192[ 9 ];
	assign fresh_wire_458[ 10 ] = fresh_wire_192[ 10 ];
	assign fresh_wire_458[ 11 ] = fresh_wire_192[ 11 ];
	assign fresh_wire_458[ 12 ] = fresh_wire_192[ 12 ];
	assign fresh_wire_458[ 13 ] = fresh_wire_192[ 13 ];
	assign fresh_wire_458[ 14 ] = fresh_wire_192[ 14 ];
	assign fresh_wire_458[ 15 ] = fresh_wire_192[ 15 ];
	assign fresh_wire_460[ 0 ] = fresh_wire_317[ 0 ];
	assign fresh_wire_461[ 0 ] = fresh_wire_459[ 0 ];
	assign fresh_wire_461[ 1 ] = fresh_wire_459[ 1 ];
	assign fresh_wire_461[ 2 ] = fresh_wire_459[ 2 ];
	assign fresh_wire_461[ 3 ] = fresh_wire_459[ 3 ];
	assign fresh_wire_461[ 4 ] = fresh_wire_459[ 4 ];
	assign fresh_wire_461[ 5 ] = fresh_wire_459[ 5 ];
	assign fresh_wire_461[ 6 ] = fresh_wire_459[ 6 ];
	assign fresh_wire_461[ 7 ] = fresh_wire_459[ 7 ];
	assign fresh_wire_461[ 8 ] = fresh_wire_459[ 8 ];
	assign fresh_wire_461[ 9 ] = fresh_wire_459[ 9 ];
	assign fresh_wire_461[ 10 ] = fresh_wire_459[ 10 ];
	assign fresh_wire_461[ 11 ] = fresh_wire_459[ 11 ];
	assign fresh_wire_461[ 12 ] = fresh_wire_459[ 12 ];
	assign fresh_wire_461[ 13 ] = fresh_wire_459[ 13 ];
	assign fresh_wire_461[ 14 ] = fresh_wire_459[ 14 ];
	assign fresh_wire_461[ 15 ] = fresh_wire_459[ 15 ];
	assign fresh_wire_462[ 0 ] = fresh_wire_604[ 0 ];
	assign fresh_wire_462[ 1 ] = fresh_wire_604[ 1 ];
	assign fresh_wire_462[ 2 ] = fresh_wire_604[ 2 ];
	assign fresh_wire_462[ 3 ] = fresh_wire_604[ 3 ];
	assign fresh_wire_462[ 4 ] = fresh_wire_604[ 4 ];
	assign fresh_wire_462[ 5 ] = fresh_wire_604[ 5 ];
	assign fresh_wire_462[ 6 ] = fresh_wire_604[ 6 ];
	assign fresh_wire_462[ 7 ] = fresh_wire_604[ 7 ];
	assign fresh_wire_462[ 8 ] = fresh_wire_604[ 8 ];
	assign fresh_wire_462[ 9 ] = fresh_wire_604[ 9 ];
	assign fresh_wire_462[ 10 ] = fresh_wire_604[ 10 ];
	assign fresh_wire_462[ 11 ] = fresh_wire_604[ 11 ];
	assign fresh_wire_462[ 12 ] = fresh_wire_604[ 12 ];
	assign fresh_wire_462[ 13 ] = fresh_wire_604[ 13 ];
	assign fresh_wire_462[ 14 ] = fresh_wire_604[ 14 ];
	assign fresh_wire_462[ 15 ] = fresh_wire_604[ 15 ];
	assign fresh_wire_464[ 0 ] = fresh_wire_310[ 0 ];
	assign fresh_wire_465[ 0 ] = fresh_wire_463[ 0 ];
	assign fresh_wire_465[ 1 ] = fresh_wire_463[ 1 ];
	assign fresh_wire_465[ 2 ] = fresh_wire_463[ 2 ];
	assign fresh_wire_465[ 3 ] = fresh_wire_463[ 3 ];
	assign fresh_wire_465[ 4 ] = fresh_wire_463[ 4 ];
	assign fresh_wire_465[ 5 ] = fresh_wire_463[ 5 ];
	assign fresh_wire_465[ 6 ] = fresh_wire_463[ 6 ];
	assign fresh_wire_465[ 7 ] = fresh_wire_463[ 7 ];
	assign fresh_wire_465[ 8 ] = fresh_wire_463[ 8 ];
	assign fresh_wire_465[ 9 ] = fresh_wire_463[ 9 ];
	assign fresh_wire_465[ 10 ] = fresh_wire_463[ 10 ];
	assign fresh_wire_465[ 11 ] = fresh_wire_463[ 11 ];
	assign fresh_wire_465[ 12 ] = fresh_wire_463[ 12 ];
	assign fresh_wire_465[ 13 ] = fresh_wire_463[ 13 ];
	assign fresh_wire_465[ 14 ] = fresh_wire_463[ 14 ];
	assign fresh_wire_465[ 15 ] = fresh_wire_463[ 15 ];
	assign fresh_wire_466[ 0 ] = fresh_wire_406[ 0 ];
	assign fresh_wire_466[ 1 ] = fresh_wire_406[ 1 ];
	assign fresh_wire_466[ 2 ] = fresh_wire_406[ 2 ];
	assign fresh_wire_466[ 3 ] = fresh_wire_406[ 3 ];
	assign fresh_wire_466[ 4 ] = fresh_wire_406[ 4 ];
	assign fresh_wire_466[ 5 ] = fresh_wire_406[ 5 ];
	assign fresh_wire_466[ 6 ] = fresh_wire_406[ 6 ];
	assign fresh_wire_466[ 7 ] = fresh_wire_406[ 7 ];
	assign fresh_wire_466[ 8 ] = fresh_wire_406[ 8 ];
	assign fresh_wire_466[ 9 ] = fresh_wire_406[ 9 ];
	assign fresh_wire_466[ 10 ] = fresh_wire_406[ 10 ];
	assign fresh_wire_466[ 11 ] = fresh_wire_406[ 11 ];
	assign fresh_wire_466[ 12 ] = fresh_wire_406[ 12 ];
	assign fresh_wire_466[ 13 ] = fresh_wire_406[ 13 ];
	assign fresh_wire_466[ 14 ] = fresh_wire_406[ 14 ];
	assign fresh_wire_466[ 15 ] = fresh_wire_406[ 15 ];
	assign fresh_wire_468[ 0 ] = fresh_wire_298[ 0 ];
	assign fresh_wire_469[ 0 ] = fresh_wire_406[ 0 ];
	assign fresh_wire_469[ 1 ] = fresh_wire_406[ 1 ];
	assign fresh_wire_469[ 2 ] = fresh_wire_406[ 2 ];
	assign fresh_wire_469[ 3 ] = fresh_wire_406[ 3 ];
	assign fresh_wire_469[ 4 ] = fresh_wire_406[ 4 ];
	assign fresh_wire_469[ 5 ] = fresh_wire_406[ 5 ];
	assign fresh_wire_469[ 6 ] = fresh_wire_406[ 6 ];
	assign fresh_wire_469[ 7 ] = fresh_wire_406[ 7 ];
	assign fresh_wire_469[ 8 ] = fresh_wire_406[ 8 ];
	assign fresh_wire_469[ 9 ] = fresh_wire_406[ 9 ];
	assign fresh_wire_469[ 10 ] = fresh_wire_406[ 10 ];
	assign fresh_wire_469[ 11 ] = fresh_wire_406[ 11 ];
	assign fresh_wire_469[ 12 ] = fresh_wire_406[ 12 ];
	assign fresh_wire_469[ 13 ] = fresh_wire_406[ 13 ];
	assign fresh_wire_469[ 14 ] = fresh_wire_406[ 14 ];
	assign fresh_wire_469[ 15 ] = fresh_wire_406[ 15 ];
	assign fresh_wire_470[ 0 ] = fresh_wire_467[ 0 ];
	assign fresh_wire_470[ 1 ] = fresh_wire_467[ 1 ];
	assign fresh_wire_470[ 2 ] = fresh_wire_467[ 2 ];
	assign fresh_wire_470[ 3 ] = fresh_wire_467[ 3 ];
	assign fresh_wire_470[ 4 ] = fresh_wire_467[ 4 ];
	assign fresh_wire_470[ 5 ] = fresh_wire_467[ 5 ];
	assign fresh_wire_470[ 6 ] = fresh_wire_467[ 6 ];
	assign fresh_wire_470[ 7 ] = fresh_wire_467[ 7 ];
	assign fresh_wire_470[ 8 ] = fresh_wire_467[ 8 ];
	assign fresh_wire_470[ 9 ] = fresh_wire_467[ 9 ];
	assign fresh_wire_470[ 10 ] = fresh_wire_467[ 10 ];
	assign fresh_wire_470[ 11 ] = fresh_wire_467[ 11 ];
	assign fresh_wire_470[ 12 ] = fresh_wire_467[ 12 ];
	assign fresh_wire_470[ 13 ] = fresh_wire_467[ 13 ];
	assign fresh_wire_470[ 14 ] = fresh_wire_467[ 14 ];
	assign fresh_wire_470[ 15 ] = fresh_wire_467[ 15 ];
	assign fresh_wire_472[ 0 ] = fresh_wire_219[ 0 ];
	assign fresh_wire_473[ 0 ] = fresh_wire_402[ 0 ];
	assign fresh_wire_473[ 1 ] = fresh_wire_402[ 1 ];
	assign fresh_wire_474[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_474[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_476[ 0 ] = fresh_wire_329[ 0 ];
	assign fresh_wire_477[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_477[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_478[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_478[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_480[ 0 ] = fresh_wire_322[ 0 ];
	assign fresh_wire_481[ 0 ] = fresh_wire_475[ 0 ];
	assign fresh_wire_481[ 1 ] = fresh_wire_475[ 1 ];
	assign fresh_wire_482[ 0 ] = fresh_wire_479[ 0 ];
	assign fresh_wire_482[ 1 ] = fresh_wire_479[ 1 ];
	assign fresh_wire_484[ 0 ] = fresh_wire_317[ 0 ];
	assign fresh_wire_485[ 0 ] = fresh_wire_483[ 0 ];
	assign fresh_wire_485[ 1 ] = fresh_wire_483[ 1 ];
	assign fresh_wire_486[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_486[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_488[ 0 ] = fresh_wire_310[ 0 ];
	assign fresh_wire_489[ 0 ] = fresh_wire_487[ 0 ];
	assign fresh_wire_489[ 1 ] = fresh_wire_487[ 1 ];
	assign fresh_wire_490[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_490[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_492[ 0 ] = fresh_wire_298[ 0 ];
	assign fresh_wire_493[ 0 ] = fresh_wire_402[ 0 ];
	assign fresh_wire_493[ 1 ] = fresh_wire_402[ 1 ];
	assign fresh_wire_494[ 0 ] = fresh_wire_491[ 0 ];
	assign fresh_wire_494[ 1 ] = fresh_wire_491[ 1 ];
	assign fresh_wire_496[ 0 ] = fresh_wire_219[ 0 ];
	assign fresh_wire_497[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_498[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_500[ 0 ] = fresh_wire_317[ 0 ];
	assign fresh_wire_501[ 0 ] = fresh_wire_499[ 0 ];
	assign fresh_wire_502[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_504[ 0 ] = fresh_wire_310[ 0 ];
	assign fresh_wire_505[ 0 ] = fresh_wire_503[ 0 ];
	assign fresh_wire_506[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_508[ 0 ] = fresh_wire_298[ 0 ];
	assign fresh_wire_509[ 0 ] = fresh_wire_398[ 0 ];
	assign fresh_wire_510[ 0 ] = fresh_wire_507[ 0 ];
	assign fresh_wire_512[ 0 ] = fresh_wire_219[ 0 ];
	assign fresh_wire_513[ 0 ] = fresh_wire_394[ 0 ];
	assign fresh_wire_514[ 0 ] = fresh_wire_370[ 0 ];
	assign fresh_wire_516[ 0 ] = fresh_wire_329[ 0 ];
	assign fresh_wire_517[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_518[ 0 ] = fresh_wire_394[ 0 ];
	assign fresh_wire_520[ 0 ] = fresh_wire_322[ 0 ];
	assign fresh_wire_521[ 0 ] = fresh_wire_515[ 0 ];
	assign fresh_wire_522[ 0 ] = fresh_wire_519[ 0 ];
	assign fresh_wire_524[ 0 ] = fresh_wire_317[ 0 ];
	assign fresh_wire_525[ 0 ] = fresh_wire_523[ 0 ];
	assign fresh_wire_526[ 0 ] = fresh_wire_394[ 0 ];
	assign fresh_wire_528[ 0 ] = fresh_wire_310[ 0 ];
	assign fresh_wire_529[ 0 ] = fresh_wire_527[ 0 ];
	assign fresh_wire_530[ 0 ] = fresh_wire_370[ 0 ];
	assign fresh_wire_532[ 0 ] = fresh_wire_298[ 0 ];
	assign fresh_wire_533[ 0 ] = fresh_wire_394[ 0 ];
	assign fresh_wire_534[ 0 ] = fresh_wire_531[ 0 ];
	assign fresh_wire_536[ 0 ] = fresh_wire_219[ 0 ];
	assign fresh_wire_537[ 0 ] = fresh_wire_418[ 0 ];
	assign fresh_wire_537[ 1 ] = fresh_wire_418[ 1 ];
	assign fresh_wire_537[ 2 ] = fresh_wire_418[ 2 ];
	assign fresh_wire_537[ 3 ] = fresh_wire_418[ 3 ];
	assign fresh_wire_537[ 4 ] = fresh_wire_418[ 4 ];
	assign fresh_wire_537[ 5 ] = fresh_wire_418[ 5 ];
	assign fresh_wire_537[ 6 ] = fresh_wire_418[ 6 ];
	assign fresh_wire_537[ 7 ] = fresh_wire_418[ 7 ];
	assign fresh_wire_537[ 8 ] = fresh_wire_418[ 8 ];
	assign fresh_wire_537[ 9 ] = fresh_wire_418[ 9 ];
	assign fresh_wire_537[ 10 ] = fresh_wire_418[ 10 ];
	assign fresh_wire_537[ 11 ] = fresh_wire_418[ 11 ];
	assign fresh_wire_537[ 12 ] = fresh_wire_418[ 12 ];
	assign fresh_wire_537[ 13 ] = fresh_wire_418[ 13 ];
	assign fresh_wire_537[ 14 ] = fresh_wire_418[ 14 ];
	assign fresh_wire_537[ 15 ] = fresh_wire_418[ 15 ];
	assign fresh_wire_538[ 0 ] = fresh_wire_597[ 0 ];
	assign fresh_wire_538[ 1 ] = fresh_wire_597[ 1 ];
	assign fresh_wire_538[ 2 ] = fresh_wire_597[ 2 ];
	assign fresh_wire_538[ 3 ] = fresh_wire_597[ 3 ];
	assign fresh_wire_538[ 4 ] = fresh_wire_597[ 4 ];
	assign fresh_wire_538[ 5 ] = fresh_wire_597[ 5 ];
	assign fresh_wire_538[ 6 ] = fresh_wire_597[ 6 ];
	assign fresh_wire_538[ 7 ] = fresh_wire_597[ 7 ];
	assign fresh_wire_538[ 8 ] = fresh_wire_597[ 8 ];
	assign fresh_wire_538[ 9 ] = fresh_wire_597[ 9 ];
	assign fresh_wire_538[ 10 ] = fresh_wire_597[ 10 ];
	assign fresh_wire_538[ 11 ] = fresh_wire_597[ 11 ];
	assign fresh_wire_538[ 12 ] = fresh_wire_597[ 12 ];
	assign fresh_wire_538[ 13 ] = fresh_wire_597[ 13 ];
	assign fresh_wire_538[ 14 ] = fresh_wire_597[ 14 ];
	assign fresh_wire_538[ 15 ] = fresh_wire_597[ 15 ];
	assign fresh_wire_540[ 0 ] = fresh_wire_228[ 0 ];
	assign fresh_wire_541[ 0 ] = fresh_wire_418[ 0 ];
	assign fresh_wire_541[ 1 ] = fresh_wire_418[ 1 ];
	assign fresh_wire_541[ 2 ] = fresh_wire_418[ 2 ];
	assign fresh_wire_541[ 3 ] = fresh_wire_418[ 3 ];
	assign fresh_wire_541[ 4 ] = fresh_wire_418[ 4 ];
	assign fresh_wire_541[ 5 ] = fresh_wire_418[ 5 ];
	assign fresh_wire_541[ 6 ] = fresh_wire_418[ 6 ];
	assign fresh_wire_541[ 7 ] = fresh_wire_418[ 7 ];
	assign fresh_wire_541[ 8 ] = fresh_wire_418[ 8 ];
	assign fresh_wire_541[ 9 ] = fresh_wire_418[ 9 ];
	assign fresh_wire_541[ 10 ] = fresh_wire_418[ 10 ];
	assign fresh_wire_541[ 11 ] = fresh_wire_418[ 11 ];
	assign fresh_wire_541[ 12 ] = fresh_wire_418[ 12 ];
	assign fresh_wire_541[ 13 ] = fresh_wire_418[ 13 ];
	assign fresh_wire_541[ 14 ] = fresh_wire_418[ 14 ];
	assign fresh_wire_541[ 15 ] = fresh_wire_418[ 15 ];
	assign fresh_wire_542[ 0 ] = fresh_wire_181[ 0 ];
	assign fresh_wire_542[ 1 ] = fresh_wire_181[ 1 ];
	assign fresh_wire_542[ 2 ] = fresh_wire_181[ 2 ];
	assign fresh_wire_542[ 3 ] = fresh_wire_181[ 3 ];
	assign fresh_wire_542[ 4 ] = fresh_wire_181[ 4 ];
	assign fresh_wire_542[ 5 ] = fresh_wire_181[ 5 ];
	assign fresh_wire_542[ 6 ] = fresh_wire_181[ 6 ];
	assign fresh_wire_542[ 7 ] = fresh_wire_181[ 7 ];
	assign fresh_wire_542[ 8 ] = fresh_wire_181[ 8 ];
	assign fresh_wire_542[ 9 ] = fresh_wire_181[ 9 ];
	assign fresh_wire_542[ 10 ] = fresh_wire_181[ 10 ];
	assign fresh_wire_542[ 11 ] = fresh_wire_181[ 11 ];
	assign fresh_wire_542[ 12 ] = fresh_wire_181[ 12 ];
	assign fresh_wire_542[ 13 ] = fresh_wire_181[ 13 ];
	assign fresh_wire_542[ 14 ] = fresh_wire_181[ 14 ];
	assign fresh_wire_542[ 15 ] = fresh_wire_181[ 15 ];
	assign fresh_wire_544[ 0 ] = fresh_wire_234[ 0 ];
	assign fresh_wire_545[ 0 ] = fresh_wire_539[ 0 ];
	assign fresh_wire_545[ 1 ] = fresh_wire_539[ 1 ];
	assign fresh_wire_545[ 2 ] = fresh_wire_539[ 2 ];
	assign fresh_wire_545[ 3 ] = fresh_wire_539[ 3 ];
	assign fresh_wire_545[ 4 ] = fresh_wire_539[ 4 ];
	assign fresh_wire_545[ 5 ] = fresh_wire_539[ 5 ];
	assign fresh_wire_545[ 6 ] = fresh_wire_539[ 6 ];
	assign fresh_wire_545[ 7 ] = fresh_wire_539[ 7 ];
	assign fresh_wire_545[ 8 ] = fresh_wire_539[ 8 ];
	assign fresh_wire_545[ 9 ] = fresh_wire_539[ 9 ];
	assign fresh_wire_545[ 10 ] = fresh_wire_539[ 10 ];
	assign fresh_wire_545[ 11 ] = fresh_wire_539[ 11 ];
	assign fresh_wire_545[ 12 ] = fresh_wire_539[ 12 ];
	assign fresh_wire_545[ 13 ] = fresh_wire_539[ 13 ];
	assign fresh_wire_545[ 14 ] = fresh_wire_539[ 14 ];
	assign fresh_wire_545[ 15 ] = fresh_wire_539[ 15 ];
	assign fresh_wire_546[ 0 ] = fresh_wire_543[ 0 ];
	assign fresh_wire_546[ 1 ] = fresh_wire_543[ 1 ];
	assign fresh_wire_546[ 2 ] = fresh_wire_543[ 2 ];
	assign fresh_wire_546[ 3 ] = fresh_wire_543[ 3 ];
	assign fresh_wire_546[ 4 ] = fresh_wire_543[ 4 ];
	assign fresh_wire_546[ 5 ] = fresh_wire_543[ 5 ];
	assign fresh_wire_546[ 6 ] = fresh_wire_543[ 6 ];
	assign fresh_wire_546[ 7 ] = fresh_wire_543[ 7 ];
	assign fresh_wire_546[ 8 ] = fresh_wire_543[ 8 ];
	assign fresh_wire_546[ 9 ] = fresh_wire_543[ 9 ];
	assign fresh_wire_546[ 10 ] = fresh_wire_543[ 10 ];
	assign fresh_wire_546[ 11 ] = fresh_wire_543[ 11 ];
	assign fresh_wire_546[ 12 ] = fresh_wire_543[ 12 ];
	assign fresh_wire_546[ 13 ] = fresh_wire_543[ 13 ];
	assign fresh_wire_546[ 14 ] = fresh_wire_543[ 14 ];
	assign fresh_wire_546[ 15 ] = fresh_wire_543[ 15 ];
	assign fresh_wire_548[ 0 ] = fresh_wire_231[ 0 ];
	assign fresh_wire_549[ 0 ] = fresh_wire_176[ 0 ];
	assign fresh_wire_549[ 1 ] = fresh_wire_176[ 1 ];
	assign fresh_wire_549[ 2 ] = fresh_wire_176[ 2 ];
	assign fresh_wire_549[ 3 ] = fresh_wire_176[ 3 ];
	assign fresh_wire_549[ 4 ] = fresh_wire_176[ 4 ];
	assign fresh_wire_549[ 5 ] = fresh_wire_176[ 5 ];
	assign fresh_wire_549[ 6 ] = fresh_wire_176[ 6 ];
	assign fresh_wire_549[ 7 ] = fresh_wire_176[ 7 ];
	assign fresh_wire_549[ 8 ] = fresh_wire_176[ 8 ];
	assign fresh_wire_549[ 9 ] = fresh_wire_176[ 9 ];
	assign fresh_wire_549[ 10 ] = fresh_wire_176[ 10 ];
	assign fresh_wire_549[ 11 ] = fresh_wire_176[ 11 ];
	assign fresh_wire_549[ 12 ] = fresh_wire_176[ 12 ];
	assign fresh_wire_549[ 13 ] = fresh_wire_176[ 13 ];
	assign fresh_wire_549[ 14 ] = fresh_wire_176[ 14 ];
	assign fresh_wire_549[ 15 ] = fresh_wire_176[ 15 ];
	assign fresh_wire_550[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_550[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_550[ 2 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_550[ 3 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_550[ 4 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_550[ 5 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_550[ 6 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_550[ 7 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_550[ 8 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_550[ 9 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_550[ 10 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_550[ 11 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_550[ 12 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_550[ 13 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_550[ 14 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_550[ 15 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_552[ 0 ] = fresh_wire_261[ 0 ];
	assign fresh_wire_553[ 0 ] = fresh_wire_414[ 0 ];
	assign fresh_wire_553[ 1 ] = fresh_wire_414[ 1 ];
	assign fresh_wire_553[ 2 ] = fresh_wire_414[ 2 ];
	assign fresh_wire_553[ 3 ] = fresh_wire_414[ 3 ];
	assign fresh_wire_553[ 4 ] = fresh_wire_414[ 4 ];
	assign fresh_wire_553[ 5 ] = fresh_wire_414[ 5 ];
	assign fresh_wire_553[ 6 ] = fresh_wire_414[ 6 ];
	assign fresh_wire_553[ 7 ] = fresh_wire_414[ 7 ];
	assign fresh_wire_553[ 8 ] = fresh_wire_414[ 8 ];
	assign fresh_wire_553[ 9 ] = fresh_wire_414[ 9 ];
	assign fresh_wire_553[ 10 ] = fresh_wire_414[ 10 ];
	assign fresh_wire_553[ 11 ] = fresh_wire_414[ 11 ];
	assign fresh_wire_553[ 12 ] = fresh_wire_414[ 12 ];
	assign fresh_wire_553[ 13 ] = fresh_wire_414[ 13 ];
	assign fresh_wire_553[ 14 ] = fresh_wire_414[ 14 ];
	assign fresh_wire_553[ 15 ] = fresh_wire_414[ 15 ];
	assign fresh_wire_554[ 0 ] = fresh_wire_551[ 0 ];
	assign fresh_wire_554[ 1 ] = fresh_wire_551[ 1 ];
	assign fresh_wire_554[ 2 ] = fresh_wire_551[ 2 ];
	assign fresh_wire_554[ 3 ] = fresh_wire_551[ 3 ];
	assign fresh_wire_554[ 4 ] = fresh_wire_551[ 4 ];
	assign fresh_wire_554[ 5 ] = fresh_wire_551[ 5 ];
	assign fresh_wire_554[ 6 ] = fresh_wire_551[ 6 ];
	assign fresh_wire_554[ 7 ] = fresh_wire_551[ 7 ];
	assign fresh_wire_554[ 8 ] = fresh_wire_551[ 8 ];
	assign fresh_wire_554[ 9 ] = fresh_wire_551[ 9 ];
	assign fresh_wire_554[ 10 ] = fresh_wire_551[ 10 ];
	assign fresh_wire_554[ 11 ] = fresh_wire_551[ 11 ];
	assign fresh_wire_554[ 12 ] = fresh_wire_551[ 12 ];
	assign fresh_wire_554[ 13 ] = fresh_wire_551[ 13 ];
	assign fresh_wire_554[ 14 ] = fresh_wire_551[ 14 ];
	assign fresh_wire_554[ 15 ] = fresh_wire_551[ 15 ];
	assign fresh_wire_556[ 0 ] = fresh_wire_234[ 0 ];
	assign fresh_wire_557[ 0 ] = fresh_wire_414[ 0 ];
	assign fresh_wire_557[ 1 ] = fresh_wire_414[ 1 ];
	assign fresh_wire_557[ 2 ] = fresh_wire_414[ 2 ];
	assign fresh_wire_557[ 3 ] = fresh_wire_414[ 3 ];
	assign fresh_wire_557[ 4 ] = fresh_wire_414[ 4 ];
	assign fresh_wire_557[ 5 ] = fresh_wire_414[ 5 ];
	assign fresh_wire_557[ 6 ] = fresh_wire_414[ 6 ];
	assign fresh_wire_557[ 7 ] = fresh_wire_414[ 7 ];
	assign fresh_wire_557[ 8 ] = fresh_wire_414[ 8 ];
	assign fresh_wire_557[ 9 ] = fresh_wire_414[ 9 ];
	assign fresh_wire_557[ 10 ] = fresh_wire_414[ 10 ];
	assign fresh_wire_557[ 11 ] = fresh_wire_414[ 11 ];
	assign fresh_wire_557[ 12 ] = fresh_wire_414[ 12 ];
	assign fresh_wire_557[ 13 ] = fresh_wire_414[ 13 ];
	assign fresh_wire_557[ 14 ] = fresh_wire_414[ 14 ];
	assign fresh_wire_557[ 15 ] = fresh_wire_414[ 15 ];
	assign fresh_wire_558[ 0 ] = fresh_wire_555[ 0 ];
	assign fresh_wire_558[ 1 ] = fresh_wire_555[ 1 ];
	assign fresh_wire_558[ 2 ] = fresh_wire_555[ 2 ];
	assign fresh_wire_558[ 3 ] = fresh_wire_555[ 3 ];
	assign fresh_wire_558[ 4 ] = fresh_wire_555[ 4 ];
	assign fresh_wire_558[ 5 ] = fresh_wire_555[ 5 ];
	assign fresh_wire_558[ 6 ] = fresh_wire_555[ 6 ];
	assign fresh_wire_558[ 7 ] = fresh_wire_555[ 7 ];
	assign fresh_wire_558[ 8 ] = fresh_wire_555[ 8 ];
	assign fresh_wire_558[ 9 ] = fresh_wire_555[ 9 ];
	assign fresh_wire_558[ 10 ] = fresh_wire_555[ 10 ];
	assign fresh_wire_558[ 11 ] = fresh_wire_555[ 11 ];
	assign fresh_wire_558[ 12 ] = fresh_wire_555[ 12 ];
	assign fresh_wire_558[ 13 ] = fresh_wire_555[ 13 ];
	assign fresh_wire_558[ 14 ] = fresh_wire_555[ 14 ];
	assign fresh_wire_558[ 15 ] = fresh_wire_555[ 15 ];
	assign fresh_wire_560[ 0 ] = fresh_wire_231[ 0 ];
	assign fresh_wire_561[ 0 ] = fresh_wire_186[ 0 ];
	assign fresh_wire_561[ 1 ] = fresh_wire_186[ 1 ];
	assign fresh_wire_561[ 2 ] = fresh_wire_186[ 2 ];
	assign fresh_wire_561[ 3 ] = fresh_wire_186[ 3 ];
	assign fresh_wire_561[ 4 ] = fresh_wire_186[ 4 ];
	assign fresh_wire_561[ 5 ] = fresh_wire_186[ 5 ];
	assign fresh_wire_561[ 6 ] = fresh_wire_186[ 6 ];
	assign fresh_wire_561[ 7 ] = fresh_wire_186[ 7 ];
	assign fresh_wire_561[ 8 ] = fresh_wire_186[ 8 ];
	assign fresh_wire_561[ 9 ] = fresh_wire_186[ 9 ];
	assign fresh_wire_561[ 10 ] = fresh_wire_186[ 10 ];
	assign fresh_wire_561[ 11 ] = fresh_wire_186[ 11 ];
	assign fresh_wire_561[ 12 ] = fresh_wire_186[ 12 ];
	assign fresh_wire_561[ 13 ] = fresh_wire_186[ 13 ];
	assign fresh_wire_561[ 14 ] = fresh_wire_186[ 14 ];
	assign fresh_wire_561[ 15 ] = fresh_wire_186[ 15 ];
	assign fresh_wire_562[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_562[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_562[ 2 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_562[ 3 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_562[ 4 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_562[ 5 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_562[ 6 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_562[ 7 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_562[ 8 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_562[ 9 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_562[ 10 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_562[ 11 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_562[ 12 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_562[ 13 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_562[ 14 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_562[ 15 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_564[ 0 ] = fresh_wire_264[ 0 ];
	assign fresh_wire_565[ 0 ] = fresh_wire_410[ 0 ];
	assign fresh_wire_565[ 1 ] = fresh_wire_410[ 1 ];
	assign fresh_wire_565[ 2 ] = fresh_wire_410[ 2 ];
	assign fresh_wire_565[ 3 ] = fresh_wire_410[ 3 ];
	assign fresh_wire_565[ 4 ] = fresh_wire_410[ 4 ];
	assign fresh_wire_565[ 5 ] = fresh_wire_410[ 5 ];
	assign fresh_wire_565[ 6 ] = fresh_wire_410[ 6 ];
	assign fresh_wire_565[ 7 ] = fresh_wire_410[ 7 ];
	assign fresh_wire_565[ 8 ] = fresh_wire_410[ 8 ];
	assign fresh_wire_565[ 9 ] = fresh_wire_410[ 9 ];
	assign fresh_wire_565[ 10 ] = fresh_wire_410[ 10 ];
	assign fresh_wire_565[ 11 ] = fresh_wire_410[ 11 ];
	assign fresh_wire_565[ 12 ] = fresh_wire_410[ 12 ];
	assign fresh_wire_565[ 13 ] = fresh_wire_410[ 13 ];
	assign fresh_wire_565[ 14 ] = fresh_wire_410[ 14 ];
	assign fresh_wire_565[ 15 ] = fresh_wire_410[ 15 ];
	assign fresh_wire_566[ 0 ] = fresh_wire_563[ 0 ];
	assign fresh_wire_566[ 1 ] = fresh_wire_563[ 1 ];
	assign fresh_wire_566[ 2 ] = fresh_wire_563[ 2 ];
	assign fresh_wire_566[ 3 ] = fresh_wire_563[ 3 ];
	assign fresh_wire_566[ 4 ] = fresh_wire_563[ 4 ];
	assign fresh_wire_566[ 5 ] = fresh_wire_563[ 5 ];
	assign fresh_wire_566[ 6 ] = fresh_wire_563[ 6 ];
	assign fresh_wire_566[ 7 ] = fresh_wire_563[ 7 ];
	assign fresh_wire_566[ 8 ] = fresh_wire_563[ 8 ];
	assign fresh_wire_566[ 9 ] = fresh_wire_563[ 9 ];
	assign fresh_wire_566[ 10 ] = fresh_wire_563[ 10 ];
	assign fresh_wire_566[ 11 ] = fresh_wire_563[ 11 ];
	assign fresh_wire_566[ 12 ] = fresh_wire_563[ 12 ];
	assign fresh_wire_566[ 13 ] = fresh_wire_563[ 13 ];
	assign fresh_wire_566[ 14 ] = fresh_wire_563[ 14 ];
	assign fresh_wire_566[ 15 ] = fresh_wire_563[ 15 ];
	assign fresh_wire_568[ 0 ] = fresh_wire_228[ 0 ];
	assign fresh_wire_569[ 0 ] = fresh_wire_567[ 0 ];
	assign fresh_wire_569[ 1 ] = fresh_wire_567[ 1 ];
	assign fresh_wire_569[ 2 ] = fresh_wire_567[ 2 ];
	assign fresh_wire_569[ 3 ] = fresh_wire_567[ 3 ];
	assign fresh_wire_569[ 4 ] = fresh_wire_567[ 4 ];
	assign fresh_wire_569[ 5 ] = fresh_wire_567[ 5 ];
	assign fresh_wire_569[ 6 ] = fresh_wire_567[ 6 ];
	assign fresh_wire_569[ 7 ] = fresh_wire_567[ 7 ];
	assign fresh_wire_569[ 8 ] = fresh_wire_567[ 8 ];
	assign fresh_wire_569[ 9 ] = fresh_wire_567[ 9 ];
	assign fresh_wire_569[ 10 ] = fresh_wire_567[ 10 ];
	assign fresh_wire_569[ 11 ] = fresh_wire_567[ 11 ];
	assign fresh_wire_569[ 12 ] = fresh_wire_567[ 12 ];
	assign fresh_wire_569[ 13 ] = fresh_wire_567[ 13 ];
	assign fresh_wire_569[ 14 ] = fresh_wire_567[ 14 ];
	assign fresh_wire_569[ 15 ] = fresh_wire_567[ 15 ];
	assign fresh_wire_570[ 0 ] = fresh_wire_410[ 0 ];
	assign fresh_wire_570[ 1 ] = fresh_wire_410[ 1 ];
	assign fresh_wire_570[ 2 ] = fresh_wire_410[ 2 ];
	assign fresh_wire_570[ 3 ] = fresh_wire_410[ 3 ];
	assign fresh_wire_570[ 4 ] = fresh_wire_410[ 4 ];
	assign fresh_wire_570[ 5 ] = fresh_wire_410[ 5 ];
	assign fresh_wire_570[ 6 ] = fresh_wire_410[ 6 ];
	assign fresh_wire_570[ 7 ] = fresh_wire_410[ 7 ];
	assign fresh_wire_570[ 8 ] = fresh_wire_410[ 8 ];
	assign fresh_wire_570[ 9 ] = fresh_wire_410[ 9 ];
	assign fresh_wire_570[ 10 ] = fresh_wire_410[ 10 ];
	assign fresh_wire_570[ 11 ] = fresh_wire_410[ 11 ];
	assign fresh_wire_570[ 12 ] = fresh_wire_410[ 12 ];
	assign fresh_wire_570[ 13 ] = fresh_wire_410[ 13 ];
	assign fresh_wire_570[ 14 ] = fresh_wire_410[ 14 ];
	assign fresh_wire_570[ 15 ] = fresh_wire_410[ 15 ];
	assign fresh_wire_572[ 0 ] = fresh_wire_231[ 0 ];
	assign fresh_wire_573[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_574[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_576[ 0 ] = fresh_wire_222[ 0 ];
	assign fresh_wire_577[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_578[ 0 ] = fresh_wire_575[ 0 ];
	assign fresh_wire_580[ 0 ] = fresh_wire_219[ 0 ];
	assign fresh_wire_581[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_582[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_584[ 0 ] = fresh_wire_225[ 0 ];
	assign fresh_wire_585[ 0 ] = fresh_wire_583[ 0 ];
	assign fresh_wire_586[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_588[ 0 ] = fresh_wire_222[ 0 ];
	assign fresh_wire_589[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_590[ 0 ] = fresh_wire_587[ 0 ];
	assign fresh_wire_592[ 0 ] = fresh_wire_219[ 0 ];
	assign fresh_wire_593[ 0 ] = fresh_wire_418[ 0 ];
	assign fresh_wire_593[ 1 ] = fresh_wire_418[ 1 ];
	assign fresh_wire_593[ 2 ] = fresh_wire_418[ 2 ];
	assign fresh_wire_593[ 3 ] = fresh_wire_418[ 3 ];
	assign fresh_wire_593[ 4 ] = fresh_wire_418[ 4 ];
	assign fresh_wire_593[ 5 ] = fresh_wire_418[ 5 ];
	assign fresh_wire_593[ 6 ] = fresh_wire_418[ 6 ];
	assign fresh_wire_593[ 7 ] = fresh_wire_418[ 7 ];
	assign fresh_wire_593[ 8 ] = fresh_wire_418[ 8 ];
	assign fresh_wire_593[ 9 ] = fresh_wire_418[ 9 ];
	assign fresh_wire_593[ 10 ] = fresh_wire_418[ 10 ];
	assign fresh_wire_593[ 11 ] = fresh_wire_418[ 11 ];
	assign fresh_wire_593[ 12 ] = fresh_wire_418[ 12 ];
	assign fresh_wire_593[ 13 ] = fresh_wire_418[ 13 ];
	assign fresh_wire_593[ 14 ] = fresh_wire_418[ 14 ];
	assign fresh_wire_593[ 15 ] = fresh_wire_418[ 15 ];
	assign fresh_wire_595[ 0 ] = fresh_wire_594[ 0 ];
	assign fresh_wire_595[ 1 ] = fresh_wire_594[ 1 ];
	assign fresh_wire_595[ 2 ] = fresh_wire_594[ 2 ];
	assign fresh_wire_595[ 3 ] = fresh_wire_594[ 3 ];
	assign fresh_wire_595[ 4 ] = fresh_wire_594[ 4 ];
	assign fresh_wire_595[ 5 ] = fresh_wire_594[ 5 ];
	assign fresh_wire_595[ 6 ] = fresh_wire_594[ 6 ];
	assign fresh_wire_595[ 7 ] = fresh_wire_594[ 7 ];
	assign fresh_wire_595[ 8 ] = fresh_wire_594[ 8 ];
	assign fresh_wire_595[ 9 ] = fresh_wire_594[ 9 ];
	assign fresh_wire_595[ 10 ] = fresh_wire_594[ 10 ];
	assign fresh_wire_595[ 11 ] = fresh_wire_594[ 11 ];
	assign fresh_wire_595[ 12 ] = fresh_wire_594[ 12 ];
	assign fresh_wire_595[ 13 ] = fresh_wire_594[ 13 ];
	assign fresh_wire_595[ 14 ] = fresh_wire_594[ 14 ];
	assign fresh_wire_595[ 15 ] = fresh_wire_594[ 15 ];
	assign fresh_wire_595[ 16 ] = fresh_wire_594[ 16 ];
	assign fresh_wire_595[ 17 ] = fresh_wire_594[ 17 ];
	assign fresh_wire_595[ 18 ] = fresh_wire_594[ 18 ];
	assign fresh_wire_595[ 19 ] = fresh_wire_594[ 19 ];
	assign fresh_wire_595[ 20 ] = fresh_wire_594[ 20 ];
	assign fresh_wire_595[ 21 ] = fresh_wire_594[ 21 ];
	assign fresh_wire_595[ 22 ] = fresh_wire_594[ 22 ];
	assign fresh_wire_595[ 23 ] = fresh_wire_594[ 23 ];
	assign fresh_wire_595[ 24 ] = fresh_wire_594[ 24 ];
	assign fresh_wire_595[ 25 ] = fresh_wire_594[ 25 ];
	assign fresh_wire_595[ 26 ] = fresh_wire_594[ 26 ];
	assign fresh_wire_595[ 27 ] = fresh_wire_594[ 27 ];
	assign fresh_wire_595[ 28 ] = fresh_wire_594[ 28 ];
	assign fresh_wire_595[ 29 ] = fresh_wire_594[ 29 ];
	assign fresh_wire_595[ 30 ] = fresh_wire_594[ 30 ];
	assign fresh_wire_595[ 31 ] = fresh_wire_594[ 31 ];
	assign fresh_wire_596[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 1 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_596[ 2 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 3 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 4 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 5 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 6 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 7 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 8 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 9 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 10 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 11 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 12 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 13 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 14 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 15 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 16 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 17 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 18 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 19 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 20 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 21 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 22 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 23 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 24 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 25 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 26 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 27 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 28 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 29 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 30 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_596[ 31 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_598[ 0 ] = fresh_wire_939[ 0 ];
	assign fresh_wire_598[ 1 ] = fresh_wire_939[ 1 ];
	assign fresh_wire_598[ 2 ] = fresh_wire_939[ 2 ];
	assign fresh_wire_598[ 3 ] = fresh_wire_939[ 3 ];
	assign fresh_wire_598[ 4 ] = fresh_wire_939[ 4 ];
	assign fresh_wire_598[ 5 ] = fresh_wire_939[ 5 ];
	assign fresh_wire_598[ 6 ] = fresh_wire_939[ 6 ];
	assign fresh_wire_598[ 7 ] = fresh_wire_939[ 7 ];
	assign fresh_wire_598[ 8 ] = fresh_wire_939[ 8 ];
	assign fresh_wire_598[ 9 ] = fresh_wire_939[ 9 ];
	assign fresh_wire_598[ 10 ] = fresh_wire_939[ 10 ];
	assign fresh_wire_598[ 11 ] = fresh_wire_939[ 11 ];
	assign fresh_wire_598[ 12 ] = fresh_wire_939[ 12 ];
	assign fresh_wire_598[ 13 ] = fresh_wire_939[ 13 ];
	assign fresh_wire_598[ 14 ] = fresh_wire_939[ 14 ];
	assign fresh_wire_598[ 15 ] = fresh_wire_939[ 15 ];
	assign fresh_wire_598[ 16 ] = fresh_wire_1037[ 0 ];
	assign fresh_wire_598[ 17 ] = fresh_wire_1037[ 1 ];
	assign fresh_wire_598[ 18 ] = fresh_wire_1037[ 2 ];
	assign fresh_wire_598[ 19 ] = fresh_wire_1037[ 3 ];
	assign fresh_wire_598[ 20 ] = fresh_wire_1037[ 4 ];
	assign fresh_wire_598[ 21 ] = fresh_wire_1037[ 5 ];
	assign fresh_wire_598[ 22 ] = fresh_wire_1037[ 6 ];
	assign fresh_wire_598[ 23 ] = fresh_wire_1037[ 7 ];
	assign fresh_wire_598[ 24 ] = fresh_wire_1037[ 8 ];
	assign fresh_wire_598[ 25 ] = fresh_wire_1037[ 9 ];
	assign fresh_wire_598[ 26 ] = fresh_wire_1037[ 10 ];
	assign fresh_wire_598[ 27 ] = fresh_wire_1037[ 11 ];
	assign fresh_wire_598[ 28 ] = fresh_wire_1037[ 12 ];
	assign fresh_wire_598[ 29 ] = fresh_wire_1037[ 13 ];
	assign fresh_wire_598[ 30 ] = fresh_wire_1037[ 14 ];
	assign fresh_wire_598[ 31 ] = fresh_wire_1037[ 15 ];
	assign fresh_wire_599[ 0 ] = fresh_wire_714[ 0 ];
	assign fresh_wire_599[ 1 ] = fresh_wire_714[ 1 ];
	assign fresh_wire_599[ 2 ] = fresh_wire_714[ 2 ];
	assign fresh_wire_599[ 3 ] = fresh_wire_714[ 3 ];
	assign fresh_wire_599[ 4 ] = fresh_wire_714[ 4 ];
	assign fresh_wire_599[ 5 ] = fresh_wire_714[ 5 ];
	assign fresh_wire_599[ 6 ] = fresh_wire_714[ 6 ];
	assign fresh_wire_599[ 7 ] = fresh_wire_714[ 7 ];
	assign fresh_wire_599[ 8 ] = fresh_wire_714[ 8 ];
	assign fresh_wire_599[ 9 ] = fresh_wire_714[ 9 ];
	assign fresh_wire_599[ 10 ] = fresh_wire_714[ 10 ];
	assign fresh_wire_599[ 11 ] = fresh_wire_714[ 11 ];
	assign fresh_wire_599[ 12 ] = fresh_wire_714[ 12 ];
	assign fresh_wire_599[ 13 ] = fresh_wire_714[ 13 ];
	assign fresh_wire_599[ 14 ] = fresh_wire_714[ 14 ];
	assign fresh_wire_599[ 15 ] = fresh_wire_714[ 15 ];
	assign fresh_wire_599[ 16 ] = fresh_wire_714[ 16 ];
	assign fresh_wire_599[ 17 ] = fresh_wire_714[ 17 ];
	assign fresh_wire_599[ 18 ] = fresh_wire_714[ 18 ];
	assign fresh_wire_599[ 19 ] = fresh_wire_714[ 19 ];
	assign fresh_wire_599[ 20 ] = fresh_wire_714[ 20 ];
	assign fresh_wire_599[ 21 ] = fresh_wire_714[ 21 ];
	assign fresh_wire_599[ 22 ] = fresh_wire_714[ 22 ];
	assign fresh_wire_599[ 23 ] = fresh_wire_714[ 23 ];
	assign fresh_wire_599[ 24 ] = fresh_wire_714[ 24 ];
	assign fresh_wire_599[ 25 ] = fresh_wire_714[ 25 ];
	assign fresh_wire_599[ 26 ] = fresh_wire_714[ 26 ];
	assign fresh_wire_599[ 27 ] = fresh_wire_714[ 27 ];
	assign fresh_wire_599[ 28 ] = fresh_wire_714[ 28 ];
	assign fresh_wire_599[ 29 ] = fresh_wire_714[ 29 ];
	assign fresh_wire_599[ 30 ] = fresh_wire_714[ 30 ];
	assign fresh_wire_599[ 31 ] = fresh_wire_714[ 31 ];
	assign fresh_wire_601[ 0 ] = fresh_wire_216[ 0 ];
	assign fresh_wire_602[ 0 ] = fresh_wire_192[ 0 ];
	assign fresh_wire_602[ 1 ] = fresh_wire_192[ 1 ];
	assign fresh_wire_602[ 2 ] = fresh_wire_192[ 2 ];
	assign fresh_wire_602[ 3 ] = fresh_wire_192[ 3 ];
	assign fresh_wire_602[ 4 ] = fresh_wire_192[ 4 ];
	assign fresh_wire_602[ 5 ] = fresh_wire_192[ 5 ];
	assign fresh_wire_602[ 6 ] = fresh_wire_192[ 6 ];
	assign fresh_wire_602[ 7 ] = fresh_wire_192[ 7 ];
	assign fresh_wire_602[ 8 ] = fresh_wire_192[ 8 ];
	assign fresh_wire_602[ 9 ] = fresh_wire_192[ 9 ];
	assign fresh_wire_602[ 10 ] = fresh_wire_192[ 10 ];
	assign fresh_wire_602[ 11 ] = fresh_wire_192[ 11 ];
	assign fresh_wire_602[ 12 ] = fresh_wire_192[ 12 ];
	assign fresh_wire_602[ 13 ] = fresh_wire_192[ 13 ];
	assign fresh_wire_602[ 14 ] = fresh_wire_192[ 14 ];
	assign fresh_wire_602[ 15 ] = fresh_wire_192[ 15 ];
	assign fresh_wire_603[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_603[ 1 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_603[ 2 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_603[ 3 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_603[ 4 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_603[ 5 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_603[ 6 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_603[ 7 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_603[ 8 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_603[ 9 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_603[ 10 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_603[ 11 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_603[ 12 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_603[ 13 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_603[ 14 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_603[ 15 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_605[ 0 ] = fresh_wire_243[ 0 ];
	assign fresh_wire_607[ 0 ] = fresh_wire_878[ 0 ];
	assign fresh_wire_607[ 1 ] = fresh_wire_878[ 1 ];
	assign fresh_wire_607[ 2 ] = fresh_wire_878[ 2 ];
	assign fresh_wire_607[ 3 ] = fresh_wire_878[ 3 ];
	assign fresh_wire_607[ 4 ] = fresh_wire_878[ 4 ];
	assign fresh_wire_607[ 5 ] = fresh_wire_878[ 5 ];
	assign fresh_wire_607[ 6 ] = fresh_wire_878[ 6 ];
	assign fresh_wire_607[ 7 ] = fresh_wire_878[ 7 ];
	assign fresh_wire_607[ 8 ] = fresh_wire_878[ 8 ];
	assign fresh_wire_607[ 9 ] = fresh_wire_878[ 9 ];
	assign fresh_wire_607[ 10 ] = fresh_wire_878[ 10 ];
	assign fresh_wire_607[ 11 ] = fresh_wire_878[ 11 ];
	assign fresh_wire_607[ 12 ] = fresh_wire_878[ 12 ];
	assign fresh_wire_607[ 13 ] = fresh_wire_878[ 13 ];
	assign fresh_wire_607[ 14 ] = fresh_wire_878[ 14 ];
	assign fresh_wire_607[ 15 ] = fresh_wire_878[ 15 ];
	assign fresh_wire_608[ 0 ] = fresh_wire_379[ 0 ];
	assign fresh_wire_608[ 1 ] = fresh_wire_379[ 1 ];
	assign fresh_wire_608[ 2 ] = fresh_wire_379[ 2 ];
	assign fresh_wire_608[ 3 ] = fresh_wire_379[ 3 ];
	assign fresh_wire_608[ 4 ] = fresh_wire_379[ 4 ];
	assign fresh_wire_608[ 5 ] = fresh_wire_379[ 5 ];
	assign fresh_wire_608[ 6 ] = fresh_wire_379[ 6 ];
	assign fresh_wire_608[ 7 ] = fresh_wire_379[ 7 ];
	assign fresh_wire_608[ 8 ] = fresh_wire_379[ 8 ];
	assign fresh_wire_608[ 9 ] = fresh_wire_379[ 9 ];
	assign fresh_wire_608[ 10 ] = fresh_wire_379[ 10 ];
	assign fresh_wire_608[ 11 ] = fresh_wire_379[ 11 ];
	assign fresh_wire_608[ 12 ] = fresh_wire_379[ 12 ];
	assign fresh_wire_608[ 13 ] = fresh_wire_379[ 13 ];
	assign fresh_wire_608[ 14 ] = fresh_wire_379[ 14 ];
	assign fresh_wire_608[ 15 ] = fresh_wire_379[ 15 ];
	assign fresh_wire_610[ 0 ] = fresh_wire_258[ 0 ];
	assign fresh_wire_611[ 0 ] = fresh_wire_666[ 0 ];
	assign fresh_wire_611[ 1 ] = fresh_wire_666[ 1 ];
	assign fresh_wire_612[ 0 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_612[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_614[ 0 ] = fresh_wire_426[ 0 ];
	assign fresh_wire_615[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_617[ 0 ] = fresh_wire_422[ 0 ];
	assign fresh_wire_618[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_620[ 0 ] = fresh_wire_426[ 0 ];
	assign fresh_wire_621[ 0 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_623[ 0 ] = fresh_wire_666[ 0 ];
	assign fresh_wire_623[ 1 ] = fresh_wire_666[ 1 ];
	assign fresh_wire_624[ 0 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_624[ 1 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_626[ 0 ] = fresh_wire_666[ 0 ];
	assign fresh_wire_626[ 1 ] = fresh_wire_666[ 1 ];
	assign fresh_wire_627[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_627[ 1 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_629[ 0 ] = fresh_wire_422[ 0 ];
	assign fresh_wire_630[ 0 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_632[ 0 ] = fresh_wire_666[ 0 ];
	assign fresh_wire_632[ 1 ] = fresh_wire_666[ 1 ];
	assign fresh_wire_633[ 0 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_633[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_635[ 0 ] = fresh_wire_666[ 0 ];
	assign fresh_wire_635[ 1 ] = fresh_wire_666[ 1 ];
	assign fresh_wire_636[ 0 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_636[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_638[ 0 ] = fresh_wire_616[ 0 ];
	assign fresh_wire_640[ 0 ] = fresh_wire_639[ 0 ];
	assign fresh_wire_641[ 0 ] = fresh_wire_644[ 0 ];
	assign fresh_wire_643[ 0 ] = fresh_wire_619[ 0 ];
	assign fresh_wire_645[ 0 ] = fresh_wire_1170[ 0 ];
	assign fresh_wire_646[ 0 ] = fresh_wire_649[ 0 ];
	assign fresh_wire_648[ 0 ] = fresh_wire_642[ 0 ];
	assign fresh_wire_650[ 0 ] = fresh_wire_1171[ 0 ];
	assign fresh_wire_651[ 0 ] = fresh_wire_654[ 0 ];
	assign fresh_wire_653[ 0 ] = fresh_wire_622[ 0 ];
	assign fresh_wire_655[ 0 ] = fresh_wire_1172[ 0 ];
	assign fresh_wire_656[ 0 ] = fresh_wire_659[ 0 ];
	assign fresh_wire_658[ 0 ] = fresh_wire_616[ 0 ];
	assign fresh_wire_660[ 0 ] = fresh_wire_1173[ 0 ];
	assign fresh_wire_661[ 0 ] = fresh_wire_664[ 0 ];
	assign fresh_wire_663[ 0 ] = fresh_wire_622[ 0 ];
	assign fresh_wire_665[ 0 ] = fresh_wire_686[ 0 ];
	assign fresh_wire_665[ 1 ] = fresh_wire_686[ 1 ];
	assign fresh_wire_667[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_668[ 0 ] = fresh_wire_1153[ 0 ];
	assign fresh_wire_669[ 0 ] = fresh_wire_96[ 0 ];
	assign fresh_wire_669[ 1 ] = fresh_wire_94[ 0 ];
	assign fresh_wire_669[ 2 ] = fresh_wire_92[ 0 ];
	assign fresh_wire_669[ 3 ] = fresh_wire_90[ 0 ];
	assign fresh_wire_669[ 4 ] = fresh_wire_88[ 0 ];
	assign fresh_wire_669[ 5 ] = fresh_wire_86[ 0 ];
	assign fresh_wire_669[ 6 ] = fresh_wire_114[ 0 ];
	assign fresh_wire_669[ 7 ] = fresh_wire_112[ 0 ];
	assign fresh_wire_669[ 8 ] = fresh_wire_110[ 0 ];
	assign fresh_wire_669[ 9 ] = fresh_wire_108[ 0 ];
	assign fresh_wire_669[ 10 ] = fresh_wire_106[ 0 ];
	assign fresh_wire_669[ 11 ] = fresh_wire_104[ 0 ];
	assign fresh_wire_669[ 12 ] = fresh_wire_102[ 0 ];
	assign fresh_wire_669[ 13 ] = fresh_wire_100[ 0 ];
	assign fresh_wire_669[ 14 ] = fresh_wire_98[ 0 ];
	assign fresh_wire_669[ 15 ] = fresh_wire_84[ 0 ];
	assign fresh_wire_669[ 16 ] = fresh_wire_670[ 0 ];
	assign fresh_wire_669[ 17 ] = fresh_wire_670[ 1 ];
	assign fresh_wire_669[ 18 ] = fresh_wire_670[ 2 ];
	assign fresh_wire_669[ 19 ] = fresh_wire_670[ 3 ];
	assign fresh_wire_669[ 20 ] = fresh_wire_670[ 4 ];
	assign fresh_wire_669[ 21 ] = fresh_wire_670[ 5 ];
	assign fresh_wire_669[ 22 ] = fresh_wire_670[ 6 ];
	assign fresh_wire_669[ 23 ] = fresh_wire_670[ 7 ];
	assign fresh_wire_669[ 24 ] = fresh_wire_670[ 8 ];
	assign fresh_wire_669[ 25 ] = fresh_wire_670[ 9 ];
	assign fresh_wire_669[ 26 ] = fresh_wire_670[ 10 ];
	assign fresh_wire_669[ 27 ] = fresh_wire_670[ 11 ];
	assign fresh_wire_669[ 28 ] = fresh_wire_670[ 12 ];
	assign fresh_wire_669[ 29 ] = fresh_wire_670[ 13 ];
	assign fresh_wire_669[ 30 ] = fresh_wire_670[ 14 ];
	assign fresh_wire_669[ 31 ] = fresh_wire_670[ 15 ];
	assign fresh_wire_669[ 32 ] = fresh_wire_670[ 16 ];
	assign fresh_wire_669[ 33 ] = fresh_wire_670[ 17 ];
	assign fresh_wire_669[ 34 ] = fresh_wire_670[ 18 ];
	assign fresh_wire_669[ 35 ] = fresh_wire_670[ 19 ];
	assign fresh_wire_669[ 36 ] = fresh_wire_670[ 20 ];
	assign fresh_wire_669[ 37 ] = fresh_wire_670[ 21 ];
	assign fresh_wire_669[ 38 ] = fresh_wire_670[ 22 ];
	assign fresh_wire_669[ 39 ] = fresh_wire_670[ 23 ];
	assign fresh_wire_669[ 40 ] = fresh_wire_670[ 24 ];
	assign fresh_wire_669[ 41 ] = fresh_wire_670[ 25 ];
	assign fresh_wire_669[ 42 ] = fresh_wire_670[ 26 ];
	assign fresh_wire_669[ 43 ] = fresh_wire_670[ 27 ];
	assign fresh_wire_669[ 44 ] = fresh_wire_670[ 28 ];
	assign fresh_wire_669[ 45 ] = fresh_wire_670[ 29 ];
	assign fresh_wire_669[ 46 ] = fresh_wire_670[ 30 ];
	assign fresh_wire_669[ 47 ] = fresh_wire_670[ 31 ];
	assign fresh_wire_671[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_672[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_673[ 0 ] = fresh_wire_625[ 0 ];
	assign fresh_wire_675[ 0 ] = fresh_wire_662[ 0 ];
	assign fresh_wire_676[ 0 ] = fresh_wire_674[ 0 ];
	assign fresh_wire_677[ 0 ] = fresh_wire_637[ 0 ];
	assign fresh_wire_679[ 0 ] = fresh_wire_657[ 0 ];
	assign fresh_wire_680[ 0 ] = fresh_wire_666[ 0 ];
	assign fresh_wire_680[ 1 ] = fresh_wire_666[ 1 ];
	assign fresh_wire_681[ 0 ] = fresh_wire_718[ 0 ];
	assign fresh_wire_681[ 1 ] = fresh_wire_718[ 1 ];
	assign fresh_wire_683[ 0 ] = fresh_wire_652[ 0 ];
	assign fresh_wire_684[ 0 ] = fresh_wire_682[ 0 ];
	assign fresh_wire_684[ 1 ] = fresh_wire_682[ 1 ];
	assign fresh_wire_685[ 0 ] = fresh_wire_613[ 0 ];
	assign fresh_wire_685[ 1 ] = fresh_wire_613[ 1 ];
	assign fresh_wire_687[ 0 ] = fresh_wire_647[ 0 ];
	assign fresh_wire_688[ 0 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 1 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 2 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 3 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 4 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 5 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 6 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 7 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 8 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 9 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 10 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 11 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 12 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 13 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 14 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 15 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 16 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 17 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 18 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 19 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 20 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 21 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 22 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 23 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 24 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 25 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 26 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 27 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 28 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 29 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 30 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 31 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_689[ 0 ] = fresh_wire_670[ 32 ];
	assign fresh_wire_689[ 1 ] = fresh_wire_670[ 33 ];
	assign fresh_wire_689[ 2 ] = fresh_wire_670[ 34 ];
	assign fresh_wire_689[ 3 ] = fresh_wire_670[ 35 ];
	assign fresh_wire_689[ 4 ] = fresh_wire_670[ 36 ];
	assign fresh_wire_689[ 5 ] = fresh_wire_670[ 37 ];
	assign fresh_wire_689[ 6 ] = fresh_wire_670[ 38 ];
	assign fresh_wire_689[ 7 ] = fresh_wire_670[ 39 ];
	assign fresh_wire_689[ 8 ] = fresh_wire_670[ 40 ];
	assign fresh_wire_689[ 9 ] = fresh_wire_670[ 41 ];
	assign fresh_wire_689[ 10 ] = fresh_wire_670[ 42 ];
	assign fresh_wire_689[ 11 ] = fresh_wire_670[ 43 ];
	assign fresh_wire_689[ 12 ] = fresh_wire_670[ 44 ];
	assign fresh_wire_689[ 13 ] = fresh_wire_670[ 45 ];
	assign fresh_wire_689[ 14 ] = fresh_wire_670[ 46 ];
	assign fresh_wire_689[ 15 ] = fresh_wire_670[ 47 ];
	assign fresh_wire_689[ 16 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_689[ 17 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_689[ 18 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_689[ 19 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_689[ 20 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_689[ 21 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_689[ 22 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_689[ 23 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_689[ 24 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_689[ 25 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_689[ 26 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_689[ 27 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_689[ 28 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_689[ 29 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_689[ 30 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_689[ 31 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_691[ 0 ] = fresh_wire_625[ 0 ];
	assign fresh_wire_692[ 0 ] = fresh_wire_690[ 0 ];
	assign fresh_wire_692[ 1 ] = fresh_wire_690[ 1 ];
	assign fresh_wire_692[ 2 ] = fresh_wire_690[ 2 ];
	assign fresh_wire_692[ 3 ] = fresh_wire_690[ 3 ];
	assign fresh_wire_692[ 4 ] = fresh_wire_690[ 4 ];
	assign fresh_wire_692[ 5 ] = fresh_wire_690[ 5 ];
	assign fresh_wire_692[ 6 ] = fresh_wire_690[ 6 ];
	assign fresh_wire_692[ 7 ] = fresh_wire_690[ 7 ];
	assign fresh_wire_692[ 8 ] = fresh_wire_690[ 8 ];
	assign fresh_wire_692[ 9 ] = fresh_wire_690[ 9 ];
	assign fresh_wire_692[ 10 ] = fresh_wire_690[ 10 ];
	assign fresh_wire_692[ 11 ] = fresh_wire_690[ 11 ];
	assign fresh_wire_692[ 12 ] = fresh_wire_690[ 12 ];
	assign fresh_wire_692[ 13 ] = fresh_wire_690[ 13 ];
	assign fresh_wire_692[ 14 ] = fresh_wire_690[ 14 ];
	assign fresh_wire_692[ 15 ] = fresh_wire_690[ 15 ];
	assign fresh_wire_692[ 16 ] = fresh_wire_690[ 16 ];
	assign fresh_wire_692[ 17 ] = fresh_wire_690[ 17 ];
	assign fresh_wire_692[ 18 ] = fresh_wire_690[ 18 ];
	assign fresh_wire_692[ 19 ] = fresh_wire_690[ 19 ];
	assign fresh_wire_692[ 20 ] = fresh_wire_690[ 20 ];
	assign fresh_wire_692[ 21 ] = fresh_wire_690[ 21 ];
	assign fresh_wire_692[ 22 ] = fresh_wire_690[ 22 ];
	assign fresh_wire_692[ 23 ] = fresh_wire_690[ 23 ];
	assign fresh_wire_692[ 24 ] = fresh_wire_690[ 24 ];
	assign fresh_wire_692[ 25 ] = fresh_wire_690[ 25 ];
	assign fresh_wire_692[ 26 ] = fresh_wire_690[ 26 ];
	assign fresh_wire_692[ 27 ] = fresh_wire_690[ 27 ];
	assign fresh_wire_692[ 28 ] = fresh_wire_690[ 28 ];
	assign fresh_wire_692[ 29 ] = fresh_wire_690[ 29 ];
	assign fresh_wire_692[ 30 ] = fresh_wire_690[ 30 ];
	assign fresh_wire_692[ 31 ] = fresh_wire_690[ 31 ];
	assign fresh_wire_693[ 0 ] = fresh_wire_670[ 16 ];
	assign fresh_wire_693[ 1 ] = fresh_wire_670[ 17 ];
	assign fresh_wire_693[ 2 ] = fresh_wire_670[ 18 ];
	assign fresh_wire_693[ 3 ] = fresh_wire_670[ 19 ];
	assign fresh_wire_693[ 4 ] = fresh_wire_670[ 20 ];
	assign fresh_wire_693[ 5 ] = fresh_wire_670[ 21 ];
	assign fresh_wire_693[ 6 ] = fresh_wire_670[ 22 ];
	assign fresh_wire_693[ 7 ] = fresh_wire_670[ 23 ];
	assign fresh_wire_693[ 8 ] = fresh_wire_670[ 24 ];
	assign fresh_wire_693[ 9 ] = fresh_wire_670[ 25 ];
	assign fresh_wire_693[ 10 ] = fresh_wire_670[ 26 ];
	assign fresh_wire_693[ 11 ] = fresh_wire_670[ 27 ];
	assign fresh_wire_693[ 12 ] = fresh_wire_670[ 28 ];
	assign fresh_wire_693[ 13 ] = fresh_wire_670[ 29 ];
	assign fresh_wire_693[ 14 ] = fresh_wire_670[ 30 ];
	assign fresh_wire_693[ 15 ] = fresh_wire_670[ 31 ];
	assign fresh_wire_693[ 16 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_693[ 17 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_693[ 18 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_693[ 19 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_693[ 20 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_693[ 21 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_693[ 22 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_693[ 23 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_693[ 24 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_693[ 25 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_693[ 26 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_693[ 27 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_693[ 28 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_693[ 29 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_693[ 30 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_693[ 31 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_695[ 0 ] = fresh_wire_628[ 0 ];
	assign fresh_wire_696[ 0 ] = fresh_wire_694[ 0 ];
	assign fresh_wire_696[ 1 ] = fresh_wire_694[ 1 ];
	assign fresh_wire_696[ 2 ] = fresh_wire_694[ 2 ];
	assign fresh_wire_696[ 3 ] = fresh_wire_694[ 3 ];
	assign fresh_wire_696[ 4 ] = fresh_wire_694[ 4 ];
	assign fresh_wire_696[ 5 ] = fresh_wire_694[ 5 ];
	assign fresh_wire_696[ 6 ] = fresh_wire_694[ 6 ];
	assign fresh_wire_696[ 7 ] = fresh_wire_694[ 7 ];
	assign fresh_wire_696[ 8 ] = fresh_wire_694[ 8 ];
	assign fresh_wire_696[ 9 ] = fresh_wire_694[ 9 ];
	assign fresh_wire_696[ 10 ] = fresh_wire_694[ 10 ];
	assign fresh_wire_696[ 11 ] = fresh_wire_694[ 11 ];
	assign fresh_wire_696[ 12 ] = fresh_wire_694[ 12 ];
	assign fresh_wire_696[ 13 ] = fresh_wire_694[ 13 ];
	assign fresh_wire_696[ 14 ] = fresh_wire_694[ 14 ];
	assign fresh_wire_696[ 15 ] = fresh_wire_694[ 15 ];
	assign fresh_wire_696[ 16 ] = fresh_wire_694[ 16 ];
	assign fresh_wire_696[ 17 ] = fresh_wire_694[ 17 ];
	assign fresh_wire_696[ 18 ] = fresh_wire_694[ 18 ];
	assign fresh_wire_696[ 19 ] = fresh_wire_694[ 19 ];
	assign fresh_wire_696[ 20 ] = fresh_wire_694[ 20 ];
	assign fresh_wire_696[ 21 ] = fresh_wire_694[ 21 ];
	assign fresh_wire_696[ 22 ] = fresh_wire_694[ 22 ];
	assign fresh_wire_696[ 23 ] = fresh_wire_694[ 23 ];
	assign fresh_wire_696[ 24 ] = fresh_wire_694[ 24 ];
	assign fresh_wire_696[ 25 ] = fresh_wire_694[ 25 ];
	assign fresh_wire_696[ 26 ] = fresh_wire_694[ 26 ];
	assign fresh_wire_696[ 27 ] = fresh_wire_694[ 27 ];
	assign fresh_wire_696[ 28 ] = fresh_wire_694[ 28 ];
	assign fresh_wire_696[ 29 ] = fresh_wire_694[ 29 ];
	assign fresh_wire_696[ 30 ] = fresh_wire_694[ 30 ];
	assign fresh_wire_696[ 31 ] = fresh_wire_694[ 31 ];
	assign fresh_wire_697[ 0 ] = fresh_wire_670[ 0 ];
	assign fresh_wire_697[ 1 ] = fresh_wire_670[ 1 ];
	assign fresh_wire_697[ 2 ] = fresh_wire_670[ 2 ];
	assign fresh_wire_697[ 3 ] = fresh_wire_670[ 3 ];
	assign fresh_wire_697[ 4 ] = fresh_wire_670[ 4 ];
	assign fresh_wire_697[ 5 ] = fresh_wire_670[ 5 ];
	assign fresh_wire_697[ 6 ] = fresh_wire_670[ 6 ];
	assign fresh_wire_697[ 7 ] = fresh_wire_670[ 7 ];
	assign fresh_wire_697[ 8 ] = fresh_wire_670[ 8 ];
	assign fresh_wire_697[ 9 ] = fresh_wire_670[ 9 ];
	assign fresh_wire_697[ 10 ] = fresh_wire_670[ 10 ];
	assign fresh_wire_697[ 11 ] = fresh_wire_670[ 11 ];
	assign fresh_wire_697[ 12 ] = fresh_wire_670[ 12 ];
	assign fresh_wire_697[ 13 ] = fresh_wire_670[ 13 ];
	assign fresh_wire_697[ 14 ] = fresh_wire_670[ 14 ];
	assign fresh_wire_697[ 15 ] = fresh_wire_670[ 15 ];
	assign fresh_wire_697[ 16 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_697[ 17 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_697[ 18 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_697[ 19 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_697[ 20 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_697[ 21 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_697[ 22 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_697[ 23 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_697[ 24 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_697[ 25 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_697[ 26 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_697[ 27 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_697[ 28 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_697[ 29 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_697[ 30 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_697[ 31 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_699[ 0 ] = fresh_wire_634[ 0 ];
	assign fresh_wire_700[ 0 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 1 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 2 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 3 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 4 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 5 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 6 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 7 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 8 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 9 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 10 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 11 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 12 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 13 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 14 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 15 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 16 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 17 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 18 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 19 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 20 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 21 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 22 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 23 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 24 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 25 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 26 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 27 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 28 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 29 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 30 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 31 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_701[ 0 ] = fresh_wire_698[ 0 ];
	assign fresh_wire_701[ 1 ] = fresh_wire_698[ 1 ];
	assign fresh_wire_701[ 2 ] = fresh_wire_698[ 2 ];
	assign fresh_wire_701[ 3 ] = fresh_wire_698[ 3 ];
	assign fresh_wire_701[ 4 ] = fresh_wire_698[ 4 ];
	assign fresh_wire_701[ 5 ] = fresh_wire_698[ 5 ];
	assign fresh_wire_701[ 6 ] = fresh_wire_698[ 6 ];
	assign fresh_wire_701[ 7 ] = fresh_wire_698[ 7 ];
	assign fresh_wire_701[ 8 ] = fresh_wire_698[ 8 ];
	assign fresh_wire_701[ 9 ] = fresh_wire_698[ 9 ];
	assign fresh_wire_701[ 10 ] = fresh_wire_698[ 10 ];
	assign fresh_wire_701[ 11 ] = fresh_wire_698[ 11 ];
	assign fresh_wire_701[ 12 ] = fresh_wire_698[ 12 ];
	assign fresh_wire_701[ 13 ] = fresh_wire_698[ 13 ];
	assign fresh_wire_701[ 14 ] = fresh_wire_698[ 14 ];
	assign fresh_wire_701[ 15 ] = fresh_wire_698[ 15 ];
	assign fresh_wire_701[ 16 ] = fresh_wire_698[ 16 ];
	assign fresh_wire_701[ 17 ] = fresh_wire_698[ 17 ];
	assign fresh_wire_701[ 18 ] = fresh_wire_698[ 18 ];
	assign fresh_wire_701[ 19 ] = fresh_wire_698[ 19 ];
	assign fresh_wire_701[ 20 ] = fresh_wire_698[ 20 ];
	assign fresh_wire_701[ 21 ] = fresh_wire_698[ 21 ];
	assign fresh_wire_701[ 22 ] = fresh_wire_698[ 22 ];
	assign fresh_wire_701[ 23 ] = fresh_wire_698[ 23 ];
	assign fresh_wire_701[ 24 ] = fresh_wire_698[ 24 ];
	assign fresh_wire_701[ 25 ] = fresh_wire_698[ 25 ];
	assign fresh_wire_701[ 26 ] = fresh_wire_698[ 26 ];
	assign fresh_wire_701[ 27 ] = fresh_wire_698[ 27 ];
	assign fresh_wire_701[ 28 ] = fresh_wire_698[ 28 ];
	assign fresh_wire_701[ 29 ] = fresh_wire_698[ 29 ];
	assign fresh_wire_701[ 30 ] = fresh_wire_698[ 30 ];
	assign fresh_wire_701[ 31 ] = fresh_wire_698[ 31 ];
	assign fresh_wire_703[ 0 ] = fresh_wire_631[ 0 ];
	assign fresh_wire_704[ 0 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 1 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 2 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 3 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 4 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 5 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 6 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 7 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 8 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 9 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 10 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 11 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 12 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 13 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 14 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 15 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 16 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 17 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 18 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 19 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 20 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 21 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 22 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 23 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 24 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 25 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 26 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 27 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 28 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 29 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 30 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 31 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_705[ 0 ] = fresh_wire_670[ 16 ];
	assign fresh_wire_705[ 1 ] = fresh_wire_670[ 17 ];
	assign fresh_wire_705[ 2 ] = fresh_wire_670[ 18 ];
	assign fresh_wire_705[ 3 ] = fresh_wire_670[ 19 ];
	assign fresh_wire_705[ 4 ] = fresh_wire_670[ 20 ];
	assign fresh_wire_705[ 5 ] = fresh_wire_670[ 21 ];
	assign fresh_wire_705[ 6 ] = fresh_wire_670[ 22 ];
	assign fresh_wire_705[ 7 ] = fresh_wire_670[ 23 ];
	assign fresh_wire_705[ 8 ] = fresh_wire_670[ 24 ];
	assign fresh_wire_705[ 9 ] = fresh_wire_670[ 25 ];
	assign fresh_wire_705[ 10 ] = fresh_wire_670[ 26 ];
	assign fresh_wire_705[ 11 ] = fresh_wire_670[ 27 ];
	assign fresh_wire_705[ 12 ] = fresh_wire_670[ 28 ];
	assign fresh_wire_705[ 13 ] = fresh_wire_670[ 29 ];
	assign fresh_wire_705[ 14 ] = fresh_wire_670[ 30 ];
	assign fresh_wire_705[ 15 ] = fresh_wire_670[ 31 ];
	assign fresh_wire_705[ 16 ] = fresh_wire_670[ 32 ];
	assign fresh_wire_705[ 17 ] = fresh_wire_670[ 33 ];
	assign fresh_wire_705[ 18 ] = fresh_wire_670[ 34 ];
	assign fresh_wire_705[ 19 ] = fresh_wire_670[ 35 ];
	assign fresh_wire_705[ 20 ] = fresh_wire_670[ 36 ];
	assign fresh_wire_705[ 21 ] = fresh_wire_670[ 37 ];
	assign fresh_wire_705[ 22 ] = fresh_wire_670[ 38 ];
	assign fresh_wire_705[ 23 ] = fresh_wire_670[ 39 ];
	assign fresh_wire_705[ 24 ] = fresh_wire_670[ 40 ];
	assign fresh_wire_705[ 25 ] = fresh_wire_670[ 41 ];
	assign fresh_wire_705[ 26 ] = fresh_wire_670[ 42 ];
	assign fresh_wire_705[ 27 ] = fresh_wire_670[ 43 ];
	assign fresh_wire_705[ 28 ] = fresh_wire_670[ 44 ];
	assign fresh_wire_705[ 29 ] = fresh_wire_670[ 45 ];
	assign fresh_wire_705[ 30 ] = fresh_wire_670[ 46 ];
	assign fresh_wire_705[ 31 ] = fresh_wire_670[ 47 ];
	assign fresh_wire_707[ 0 ] = fresh_wire_625[ 0 ];
	assign fresh_wire_708[ 0 ] = fresh_wire_706[ 0 ];
	assign fresh_wire_708[ 1 ] = fresh_wire_706[ 1 ];
	assign fresh_wire_708[ 2 ] = fresh_wire_706[ 2 ];
	assign fresh_wire_708[ 3 ] = fresh_wire_706[ 3 ];
	assign fresh_wire_708[ 4 ] = fresh_wire_706[ 4 ];
	assign fresh_wire_708[ 5 ] = fresh_wire_706[ 5 ];
	assign fresh_wire_708[ 6 ] = fresh_wire_706[ 6 ];
	assign fresh_wire_708[ 7 ] = fresh_wire_706[ 7 ];
	assign fresh_wire_708[ 8 ] = fresh_wire_706[ 8 ];
	assign fresh_wire_708[ 9 ] = fresh_wire_706[ 9 ];
	assign fresh_wire_708[ 10 ] = fresh_wire_706[ 10 ];
	assign fresh_wire_708[ 11 ] = fresh_wire_706[ 11 ];
	assign fresh_wire_708[ 12 ] = fresh_wire_706[ 12 ];
	assign fresh_wire_708[ 13 ] = fresh_wire_706[ 13 ];
	assign fresh_wire_708[ 14 ] = fresh_wire_706[ 14 ];
	assign fresh_wire_708[ 15 ] = fresh_wire_706[ 15 ];
	assign fresh_wire_708[ 16 ] = fresh_wire_706[ 16 ];
	assign fresh_wire_708[ 17 ] = fresh_wire_706[ 17 ];
	assign fresh_wire_708[ 18 ] = fresh_wire_706[ 18 ];
	assign fresh_wire_708[ 19 ] = fresh_wire_706[ 19 ];
	assign fresh_wire_708[ 20 ] = fresh_wire_706[ 20 ];
	assign fresh_wire_708[ 21 ] = fresh_wire_706[ 21 ];
	assign fresh_wire_708[ 22 ] = fresh_wire_706[ 22 ];
	assign fresh_wire_708[ 23 ] = fresh_wire_706[ 23 ];
	assign fresh_wire_708[ 24 ] = fresh_wire_706[ 24 ];
	assign fresh_wire_708[ 25 ] = fresh_wire_706[ 25 ];
	assign fresh_wire_708[ 26 ] = fresh_wire_706[ 26 ];
	assign fresh_wire_708[ 27 ] = fresh_wire_706[ 27 ];
	assign fresh_wire_708[ 28 ] = fresh_wire_706[ 28 ];
	assign fresh_wire_708[ 29 ] = fresh_wire_706[ 29 ];
	assign fresh_wire_708[ 30 ] = fresh_wire_706[ 30 ];
	assign fresh_wire_708[ 31 ] = fresh_wire_706[ 31 ];
	assign fresh_wire_709[ 0 ] = fresh_wire_670[ 0 ];
	assign fresh_wire_709[ 1 ] = fresh_wire_670[ 1 ];
	assign fresh_wire_709[ 2 ] = fresh_wire_670[ 2 ];
	assign fresh_wire_709[ 3 ] = fresh_wire_670[ 3 ];
	assign fresh_wire_709[ 4 ] = fresh_wire_670[ 4 ];
	assign fresh_wire_709[ 5 ] = fresh_wire_670[ 5 ];
	assign fresh_wire_709[ 6 ] = fresh_wire_670[ 6 ];
	assign fresh_wire_709[ 7 ] = fresh_wire_670[ 7 ];
	assign fresh_wire_709[ 8 ] = fresh_wire_670[ 8 ];
	assign fresh_wire_709[ 9 ] = fresh_wire_670[ 9 ];
	assign fresh_wire_709[ 10 ] = fresh_wire_670[ 10 ];
	assign fresh_wire_709[ 11 ] = fresh_wire_670[ 11 ];
	assign fresh_wire_709[ 12 ] = fresh_wire_670[ 12 ];
	assign fresh_wire_709[ 13 ] = fresh_wire_670[ 13 ];
	assign fresh_wire_709[ 14 ] = fresh_wire_670[ 14 ];
	assign fresh_wire_709[ 15 ] = fresh_wire_670[ 15 ];
	assign fresh_wire_709[ 16 ] = fresh_wire_670[ 16 ];
	assign fresh_wire_709[ 17 ] = fresh_wire_670[ 17 ];
	assign fresh_wire_709[ 18 ] = fresh_wire_670[ 18 ];
	assign fresh_wire_709[ 19 ] = fresh_wire_670[ 19 ];
	assign fresh_wire_709[ 20 ] = fresh_wire_670[ 20 ];
	assign fresh_wire_709[ 21 ] = fresh_wire_670[ 21 ];
	assign fresh_wire_709[ 22 ] = fresh_wire_670[ 22 ];
	assign fresh_wire_709[ 23 ] = fresh_wire_670[ 23 ];
	assign fresh_wire_709[ 24 ] = fresh_wire_670[ 24 ];
	assign fresh_wire_709[ 25 ] = fresh_wire_670[ 25 ];
	assign fresh_wire_709[ 26 ] = fresh_wire_670[ 26 ];
	assign fresh_wire_709[ 27 ] = fresh_wire_670[ 27 ];
	assign fresh_wire_709[ 28 ] = fresh_wire_670[ 28 ];
	assign fresh_wire_709[ 29 ] = fresh_wire_670[ 29 ];
	assign fresh_wire_709[ 30 ] = fresh_wire_670[ 30 ];
	assign fresh_wire_709[ 31 ] = fresh_wire_670[ 31 ];
	assign fresh_wire_711[ 0 ] = fresh_wire_628[ 0 ];
	assign fresh_wire_712[ 0 ] = fresh_wire_702[ 0 ];
	assign fresh_wire_712[ 1 ] = fresh_wire_702[ 1 ];
	assign fresh_wire_712[ 2 ] = fresh_wire_702[ 2 ];
	assign fresh_wire_712[ 3 ] = fresh_wire_702[ 3 ];
	assign fresh_wire_712[ 4 ] = fresh_wire_702[ 4 ];
	assign fresh_wire_712[ 5 ] = fresh_wire_702[ 5 ];
	assign fresh_wire_712[ 6 ] = fresh_wire_702[ 6 ];
	assign fresh_wire_712[ 7 ] = fresh_wire_702[ 7 ];
	assign fresh_wire_712[ 8 ] = fresh_wire_702[ 8 ];
	assign fresh_wire_712[ 9 ] = fresh_wire_702[ 9 ];
	assign fresh_wire_712[ 10 ] = fresh_wire_702[ 10 ];
	assign fresh_wire_712[ 11 ] = fresh_wire_702[ 11 ];
	assign fresh_wire_712[ 12 ] = fresh_wire_702[ 12 ];
	assign fresh_wire_712[ 13 ] = fresh_wire_702[ 13 ];
	assign fresh_wire_712[ 14 ] = fresh_wire_702[ 14 ];
	assign fresh_wire_712[ 15 ] = fresh_wire_702[ 15 ];
	assign fresh_wire_712[ 16 ] = fresh_wire_702[ 16 ];
	assign fresh_wire_712[ 17 ] = fresh_wire_702[ 17 ];
	assign fresh_wire_712[ 18 ] = fresh_wire_702[ 18 ];
	assign fresh_wire_712[ 19 ] = fresh_wire_702[ 19 ];
	assign fresh_wire_712[ 20 ] = fresh_wire_702[ 20 ];
	assign fresh_wire_712[ 21 ] = fresh_wire_702[ 21 ];
	assign fresh_wire_712[ 22 ] = fresh_wire_702[ 22 ];
	assign fresh_wire_712[ 23 ] = fresh_wire_702[ 23 ];
	assign fresh_wire_712[ 24 ] = fresh_wire_702[ 24 ];
	assign fresh_wire_712[ 25 ] = fresh_wire_702[ 25 ];
	assign fresh_wire_712[ 26 ] = fresh_wire_702[ 26 ];
	assign fresh_wire_712[ 27 ] = fresh_wire_702[ 27 ];
	assign fresh_wire_712[ 28 ] = fresh_wire_702[ 28 ];
	assign fresh_wire_712[ 29 ] = fresh_wire_702[ 29 ];
	assign fresh_wire_712[ 30 ] = fresh_wire_702[ 30 ];
	assign fresh_wire_712[ 31 ] = fresh_wire_702[ 31 ];
	assign fresh_wire_713[ 0 ] = fresh_wire_710[ 0 ];
	assign fresh_wire_713[ 1 ] = fresh_wire_710[ 1 ];
	assign fresh_wire_713[ 2 ] = fresh_wire_710[ 2 ];
	assign fresh_wire_713[ 3 ] = fresh_wire_710[ 3 ];
	assign fresh_wire_713[ 4 ] = fresh_wire_710[ 4 ];
	assign fresh_wire_713[ 5 ] = fresh_wire_710[ 5 ];
	assign fresh_wire_713[ 6 ] = fresh_wire_710[ 6 ];
	assign fresh_wire_713[ 7 ] = fresh_wire_710[ 7 ];
	assign fresh_wire_713[ 8 ] = fresh_wire_710[ 8 ];
	assign fresh_wire_713[ 9 ] = fresh_wire_710[ 9 ];
	assign fresh_wire_713[ 10 ] = fresh_wire_710[ 10 ];
	assign fresh_wire_713[ 11 ] = fresh_wire_710[ 11 ];
	assign fresh_wire_713[ 12 ] = fresh_wire_710[ 12 ];
	assign fresh_wire_713[ 13 ] = fresh_wire_710[ 13 ];
	assign fresh_wire_713[ 14 ] = fresh_wire_710[ 14 ];
	assign fresh_wire_713[ 15 ] = fresh_wire_710[ 15 ];
	assign fresh_wire_713[ 16 ] = fresh_wire_710[ 16 ];
	assign fresh_wire_713[ 17 ] = fresh_wire_710[ 17 ];
	assign fresh_wire_713[ 18 ] = fresh_wire_710[ 18 ];
	assign fresh_wire_713[ 19 ] = fresh_wire_710[ 19 ];
	assign fresh_wire_713[ 20 ] = fresh_wire_710[ 20 ];
	assign fresh_wire_713[ 21 ] = fresh_wire_710[ 21 ];
	assign fresh_wire_713[ 22 ] = fresh_wire_710[ 22 ];
	assign fresh_wire_713[ 23 ] = fresh_wire_710[ 23 ];
	assign fresh_wire_713[ 24 ] = fresh_wire_710[ 24 ];
	assign fresh_wire_713[ 25 ] = fresh_wire_710[ 25 ];
	assign fresh_wire_713[ 26 ] = fresh_wire_710[ 26 ];
	assign fresh_wire_713[ 27 ] = fresh_wire_710[ 27 ];
	assign fresh_wire_713[ 28 ] = fresh_wire_710[ 28 ];
	assign fresh_wire_713[ 29 ] = fresh_wire_710[ 29 ];
	assign fresh_wire_713[ 30 ] = fresh_wire_710[ 30 ];
	assign fresh_wire_713[ 31 ] = fresh_wire_710[ 31 ];
	assign fresh_wire_715[ 0 ] = fresh_wire_622[ 0 ];
	assign fresh_wire_716[ 0 ] = fresh_wire_666[ 0 ];
	assign fresh_wire_716[ 1 ] = fresh_wire_666[ 1 ];
	assign fresh_wire_717[ 0 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_717[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_720[ 0 ] = fresh_wire_858[ 0 ];
	assign fresh_wire_720[ 1 ] = fresh_wire_858[ 1 ];
	assign fresh_wire_721[ 0 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_721[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_723[ 0 ] = fresh_wire_858[ 0 ];
	assign fresh_wire_723[ 1 ] = fresh_wire_858[ 1 ];
	assign fresh_wire_724[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_724[ 1 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_726[ 0 ] = fresh_wire_386[ 0 ];
	assign fresh_wire_727[ 0 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_729[ 0 ] = fresh_wire_382[ 0 ];
	assign fresh_wire_730[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_732[ 0 ] = fresh_wire_390[ 0 ];
	assign fresh_wire_733[ 0 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_735[ 0 ] = fresh_wire_382[ 0 ];
	assign fresh_wire_736[ 0 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_738[ 0 ] = fresh_wire_386[ 0 ];
	assign fresh_wire_739[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_741[ 0 ] = fresh_wire_390[ 0 ];
	assign fresh_wire_742[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_744[ 0 ] = fresh_wire_858[ 0 ];
	assign fresh_wire_744[ 1 ] = fresh_wire_858[ 1 ];
	assign fresh_wire_745[ 0 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_745[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_747[ 0 ] = fresh_wire_858[ 0 ];
	assign fresh_wire_747[ 1 ] = fresh_wire_858[ 1 ];
	assign fresh_wire_748[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_748[ 1 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_750[ 0 ] = fresh_wire_858[ 0 ];
	assign fresh_wire_750[ 1 ] = fresh_wire_858[ 1 ];
	assign fresh_wire_751[ 0 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_751[ 1 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_753[ 0 ] = fresh_wire_858[ 0 ];
	assign fresh_wire_753[ 1 ] = fresh_wire_858[ 1 ];
	assign fresh_wire_754[ 0 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_754[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_756[ 0 ] = fresh_wire_858[ 0 ];
	assign fresh_wire_756[ 1 ] = fresh_wire_858[ 1 ];
	assign fresh_wire_757[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_757[ 1 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_759[ 0 ] = fresh_wire_728[ 0 ];
	assign fresh_wire_761[ 0 ] = fresh_wire_760[ 0 ];
	assign fresh_wire_762[ 0 ] = fresh_wire_765[ 0 ];
	assign fresh_wire_764[ 0 ] = fresh_wire_731[ 0 ];
	assign fresh_wire_766[ 0 ] = fresh_wire_734[ 0 ];
	assign fresh_wire_768[ 0 ] = fresh_wire_767[ 0 ];
	assign fresh_wire_769[ 0 ] = fresh_wire_772[ 0 ];
	assign fresh_wire_771[ 0 ] = fresh_wire_731[ 0 ];
	assign fresh_wire_773[ 0 ] = fresh_wire_728[ 0 ];
	assign fresh_wire_775[ 0 ] = fresh_wire_774[ 0 ];
	assign fresh_wire_776[ 0 ] = fresh_wire_779[ 0 ];
	assign fresh_wire_778[ 0 ] = fresh_wire_737[ 0 ];
	assign fresh_wire_780[ 0 ] = fresh_wire_734[ 0 ];
	assign fresh_wire_782[ 0 ] = fresh_wire_781[ 0 ];
	assign fresh_wire_783[ 0 ] = fresh_wire_786[ 0 ];
	assign fresh_wire_785[ 0 ] = fresh_wire_737[ 0 ];
	assign fresh_wire_787[ 0 ] = fresh_wire_740[ 0 ];
	assign fresh_wire_789[ 0 ] = fresh_wire_788[ 0 ];
	assign fresh_wire_790[ 0 ] = fresh_wire_793[ 0 ];
	assign fresh_wire_792[ 0 ] = fresh_wire_743[ 0 ];
	assign fresh_wire_794[ 0 ] = fresh_wire_791[ 0 ];
	assign fresh_wire_796[ 0 ] = fresh_wire_795[ 0 ];
	assign fresh_wire_797[ 0 ] = fresh_wire_800[ 0 ];
	assign fresh_wire_799[ 0 ] = fresh_wire_731[ 0 ];
	assign fresh_wire_801[ 0 ] = fresh_wire_740[ 0 ];
	assign fresh_wire_803[ 0 ] = fresh_wire_802[ 0 ];
	assign fresh_wire_804[ 0 ] = fresh_wire_807[ 0 ];
	assign fresh_wire_806[ 0 ] = fresh_wire_743[ 0 ];
	assign fresh_wire_808[ 0 ] = fresh_wire_805[ 0 ];
	assign fresh_wire_810[ 0 ] = fresh_wire_809[ 0 ];
	assign fresh_wire_811[ 0 ] = fresh_wire_814[ 0 ];
	assign fresh_wire_813[ 0 ] = fresh_wire_737[ 0 ];
	assign fresh_wire_815[ 0 ] = fresh_wire_849[ 0 ];
	assign fresh_wire_817[ 0 ] = fresh_wire_816[ 0 ];
	assign fresh_wire_818[ 0 ] = fresh_wire_821[ 0 ];
	assign fresh_wire_820[ 0 ] = fresh_wire_731[ 0 ];
	assign fresh_wire_822[ 0 ] = fresh_wire_856[ 0 ];
	assign fresh_wire_824[ 0 ] = fresh_wire_823[ 0 ];
	assign fresh_wire_825[ 0 ] = fresh_wire_828[ 0 ];
	assign fresh_wire_827[ 0 ] = fresh_wire_737[ 0 ];
	assign fresh_wire_829[ 0 ] = fresh_wire_740[ 0 ];
	assign fresh_wire_831[ 0 ] = fresh_wire_830[ 0 ];
	assign fresh_wire_832[ 0 ] = fresh_wire_835[ 0 ];
	assign fresh_wire_834[ 0 ] = fresh_wire_743[ 0 ];
	assign fresh_wire_836[ 0 ] = fresh_wire_833[ 0 ];
	assign fresh_wire_838[ 0 ] = fresh_wire_837[ 0 ];
	assign fresh_wire_839[ 0 ] = fresh_wire_842[ 0 ];
	assign fresh_wire_841[ 0 ] = fresh_wire_737[ 0 ];
	assign fresh_wire_843[ 0 ] = fresh_wire_728[ 0 ];
	assign fresh_wire_845[ 0 ] = fresh_wire_734[ 0 ];
	assign fresh_wire_847[ 0 ] = fresh_wire_844[ 0 ];
	assign fresh_wire_848[ 0 ] = fresh_wire_846[ 0 ];
	assign fresh_wire_850[ 0 ] = fresh_wire_728[ 0 ];
	assign fresh_wire_852[ 0 ] = fresh_wire_734[ 0 ];
	assign fresh_wire_854[ 0 ] = fresh_wire_851[ 0 ];
	assign fresh_wire_855[ 0 ] = fresh_wire_853[ 0 ];
	assign fresh_wire_857[ 0 ] = fresh_wire_914[ 0 ];
	assign fresh_wire_857[ 1 ] = fresh_wire_914[ 1 ];
	assign fresh_wire_859[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_860[ 0 ] = fresh_wire_1153[ 0 ];
	assign fresh_wire_861[ 0 ] = fresh_wire_922[ 0 ];
	assign fresh_wire_861[ 1 ] = fresh_wire_922[ 1 ];
	assign fresh_wire_861[ 2 ] = fresh_wire_922[ 2 ];
	assign fresh_wire_861[ 3 ] = fresh_wire_922[ 3 ];
	assign fresh_wire_861[ 4 ] = fresh_wire_922[ 4 ];
	assign fresh_wire_861[ 5 ] = fresh_wire_922[ 5 ];
	assign fresh_wire_861[ 6 ] = fresh_wire_922[ 6 ];
	assign fresh_wire_861[ 7 ] = fresh_wire_922[ 7 ];
	assign fresh_wire_861[ 8 ] = fresh_wire_922[ 8 ];
	assign fresh_wire_861[ 9 ] = fresh_wire_922[ 9 ];
	assign fresh_wire_861[ 10 ] = fresh_wire_922[ 10 ];
	assign fresh_wire_861[ 11 ] = fresh_wire_922[ 11 ];
	assign fresh_wire_861[ 12 ] = fresh_wire_922[ 12 ];
	assign fresh_wire_861[ 13 ] = fresh_wire_922[ 13 ];
	assign fresh_wire_861[ 14 ] = fresh_wire_922[ 14 ];
	assign fresh_wire_861[ 15 ] = fresh_wire_922[ 15 ];
	assign fresh_wire_861[ 16 ] = fresh_wire_922[ 16 ];
	assign fresh_wire_861[ 17 ] = fresh_wire_922[ 17 ];
	assign fresh_wire_861[ 18 ] = fresh_wire_922[ 18 ];
	assign fresh_wire_861[ 19 ] = fresh_wire_922[ 19 ];
	assign fresh_wire_861[ 20 ] = fresh_wire_922[ 20 ];
	assign fresh_wire_861[ 21 ] = fresh_wire_922[ 21 ];
	assign fresh_wire_861[ 22 ] = fresh_wire_922[ 22 ];
	assign fresh_wire_861[ 23 ] = fresh_wire_922[ 23 ];
	assign fresh_wire_861[ 24 ] = fresh_wire_922[ 24 ];
	assign fresh_wire_861[ 25 ] = fresh_wire_922[ 25 ];
	assign fresh_wire_861[ 26 ] = fresh_wire_922[ 26 ];
	assign fresh_wire_861[ 27 ] = fresh_wire_922[ 27 ];
	assign fresh_wire_861[ 28 ] = fresh_wire_922[ 28 ];
	assign fresh_wire_861[ 29 ] = fresh_wire_922[ 29 ];
	assign fresh_wire_861[ 30 ] = fresh_wire_922[ 30 ];
	assign fresh_wire_861[ 31 ] = fresh_wire_922[ 31 ];
	assign fresh_wire_861[ 32 ] = fresh_wire_922[ 32 ];
	assign fresh_wire_861[ 33 ] = fresh_wire_922[ 33 ];
	assign fresh_wire_861[ 34 ] = fresh_wire_922[ 34 ];
	assign fresh_wire_861[ 35 ] = fresh_wire_922[ 35 ];
	assign fresh_wire_861[ 36 ] = fresh_wire_922[ 36 ];
	assign fresh_wire_861[ 37 ] = fresh_wire_922[ 37 ];
	assign fresh_wire_861[ 38 ] = fresh_wire_922[ 38 ];
	assign fresh_wire_861[ 39 ] = fresh_wire_922[ 39 ];
	assign fresh_wire_861[ 40 ] = fresh_wire_922[ 40 ];
	assign fresh_wire_861[ 41 ] = fresh_wire_922[ 41 ];
	assign fresh_wire_861[ 42 ] = fresh_wire_922[ 42 ];
	assign fresh_wire_861[ 43 ] = fresh_wire_922[ 43 ];
	assign fresh_wire_861[ 44 ] = fresh_wire_922[ 44 ];
	assign fresh_wire_861[ 45 ] = fresh_wire_922[ 45 ];
	assign fresh_wire_861[ 46 ] = fresh_wire_922[ 46 ];
	assign fresh_wire_861[ 47 ] = fresh_wire_922[ 47 ];
	assign fresh_wire_863[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_864[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_864[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_864[ 2 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_864[ 3 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_864[ 4 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_864[ 5 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_864[ 6 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_864[ 7 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_864[ 8 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_864[ 9 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_864[ 10 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_864[ 11 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_864[ 12 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_864[ 13 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_864[ 14 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_864[ 15 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_865[ 0 ] = fresh_wire_862[ 32 ];
	assign fresh_wire_865[ 1 ] = fresh_wire_862[ 33 ];
	assign fresh_wire_865[ 2 ] = fresh_wire_862[ 34 ];
	assign fresh_wire_865[ 3 ] = fresh_wire_862[ 35 ];
	assign fresh_wire_865[ 4 ] = fresh_wire_862[ 36 ];
	assign fresh_wire_865[ 5 ] = fresh_wire_862[ 37 ];
	assign fresh_wire_865[ 6 ] = fresh_wire_862[ 38 ];
	assign fresh_wire_865[ 7 ] = fresh_wire_862[ 39 ];
	assign fresh_wire_865[ 8 ] = fresh_wire_862[ 40 ];
	assign fresh_wire_865[ 9 ] = fresh_wire_862[ 41 ];
	assign fresh_wire_865[ 10 ] = fresh_wire_862[ 42 ];
	assign fresh_wire_865[ 11 ] = fresh_wire_862[ 43 ];
	assign fresh_wire_865[ 12 ] = fresh_wire_862[ 44 ];
	assign fresh_wire_865[ 13 ] = fresh_wire_862[ 45 ];
	assign fresh_wire_865[ 14 ] = fresh_wire_862[ 46 ];
	assign fresh_wire_865[ 15 ] = fresh_wire_862[ 47 ];
	assign fresh_wire_867[ 0 ] = fresh_wire_752[ 0 ];
	assign fresh_wire_868[ 0 ] = fresh_wire_866[ 0 ];
	assign fresh_wire_868[ 1 ] = fresh_wire_866[ 1 ];
	assign fresh_wire_868[ 2 ] = fresh_wire_866[ 2 ];
	assign fresh_wire_868[ 3 ] = fresh_wire_866[ 3 ];
	assign fresh_wire_868[ 4 ] = fresh_wire_866[ 4 ];
	assign fresh_wire_868[ 5 ] = fresh_wire_866[ 5 ];
	assign fresh_wire_868[ 6 ] = fresh_wire_866[ 6 ];
	assign fresh_wire_868[ 7 ] = fresh_wire_866[ 7 ];
	assign fresh_wire_868[ 8 ] = fresh_wire_866[ 8 ];
	assign fresh_wire_868[ 9 ] = fresh_wire_866[ 9 ];
	assign fresh_wire_868[ 10 ] = fresh_wire_866[ 10 ];
	assign fresh_wire_868[ 11 ] = fresh_wire_866[ 11 ];
	assign fresh_wire_868[ 12 ] = fresh_wire_866[ 12 ];
	assign fresh_wire_868[ 13 ] = fresh_wire_866[ 13 ];
	assign fresh_wire_868[ 14 ] = fresh_wire_866[ 14 ];
	assign fresh_wire_868[ 15 ] = fresh_wire_866[ 15 ];
	assign fresh_wire_869[ 0 ] = fresh_wire_862[ 16 ];
	assign fresh_wire_869[ 1 ] = fresh_wire_862[ 17 ];
	assign fresh_wire_869[ 2 ] = fresh_wire_862[ 18 ];
	assign fresh_wire_869[ 3 ] = fresh_wire_862[ 19 ];
	assign fresh_wire_869[ 4 ] = fresh_wire_862[ 20 ];
	assign fresh_wire_869[ 5 ] = fresh_wire_862[ 21 ];
	assign fresh_wire_869[ 6 ] = fresh_wire_862[ 22 ];
	assign fresh_wire_869[ 7 ] = fresh_wire_862[ 23 ];
	assign fresh_wire_869[ 8 ] = fresh_wire_862[ 24 ];
	assign fresh_wire_869[ 9 ] = fresh_wire_862[ 25 ];
	assign fresh_wire_869[ 10 ] = fresh_wire_862[ 26 ];
	assign fresh_wire_869[ 11 ] = fresh_wire_862[ 27 ];
	assign fresh_wire_869[ 12 ] = fresh_wire_862[ 28 ];
	assign fresh_wire_869[ 13 ] = fresh_wire_862[ 29 ];
	assign fresh_wire_869[ 14 ] = fresh_wire_862[ 30 ];
	assign fresh_wire_869[ 15 ] = fresh_wire_862[ 31 ];
	assign fresh_wire_871[ 0 ] = fresh_wire_749[ 0 ];
	assign fresh_wire_872[ 0 ] = fresh_wire_870[ 0 ];
	assign fresh_wire_872[ 1 ] = fresh_wire_870[ 1 ];
	assign fresh_wire_872[ 2 ] = fresh_wire_870[ 2 ];
	assign fresh_wire_872[ 3 ] = fresh_wire_870[ 3 ];
	assign fresh_wire_872[ 4 ] = fresh_wire_870[ 4 ];
	assign fresh_wire_872[ 5 ] = fresh_wire_870[ 5 ];
	assign fresh_wire_872[ 6 ] = fresh_wire_870[ 6 ];
	assign fresh_wire_872[ 7 ] = fresh_wire_870[ 7 ];
	assign fresh_wire_872[ 8 ] = fresh_wire_870[ 8 ];
	assign fresh_wire_872[ 9 ] = fresh_wire_870[ 9 ];
	assign fresh_wire_872[ 10 ] = fresh_wire_870[ 10 ];
	assign fresh_wire_872[ 11 ] = fresh_wire_870[ 11 ];
	assign fresh_wire_872[ 12 ] = fresh_wire_870[ 12 ];
	assign fresh_wire_872[ 13 ] = fresh_wire_870[ 13 ];
	assign fresh_wire_872[ 14 ] = fresh_wire_870[ 14 ];
	assign fresh_wire_872[ 15 ] = fresh_wire_870[ 15 ];
	assign fresh_wire_873[ 0 ] = fresh_wire_862[ 0 ];
	assign fresh_wire_873[ 1 ] = fresh_wire_862[ 1 ];
	assign fresh_wire_873[ 2 ] = fresh_wire_862[ 2 ];
	assign fresh_wire_873[ 3 ] = fresh_wire_862[ 3 ];
	assign fresh_wire_873[ 4 ] = fresh_wire_862[ 4 ];
	assign fresh_wire_873[ 5 ] = fresh_wire_862[ 5 ];
	assign fresh_wire_873[ 6 ] = fresh_wire_862[ 6 ];
	assign fresh_wire_873[ 7 ] = fresh_wire_862[ 7 ];
	assign fresh_wire_873[ 8 ] = fresh_wire_862[ 8 ];
	assign fresh_wire_873[ 9 ] = fresh_wire_862[ 9 ];
	assign fresh_wire_873[ 10 ] = fresh_wire_862[ 10 ];
	assign fresh_wire_873[ 11 ] = fresh_wire_862[ 11 ];
	assign fresh_wire_873[ 12 ] = fresh_wire_862[ 12 ];
	assign fresh_wire_873[ 13 ] = fresh_wire_862[ 13 ];
	assign fresh_wire_873[ 14 ] = fresh_wire_862[ 14 ];
	assign fresh_wire_873[ 15 ] = fresh_wire_862[ 15 ];
	assign fresh_wire_875[ 0 ] = fresh_wire_746[ 0 ];
	assign fresh_wire_876[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_876[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_876[ 2 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_876[ 3 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_876[ 4 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_876[ 5 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_876[ 6 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_876[ 7 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_876[ 8 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_876[ 9 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_876[ 10 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_876[ 11 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_876[ 12 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_876[ 13 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_876[ 14 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_876[ 15 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_877[ 0 ] = fresh_wire_874[ 0 ];
	assign fresh_wire_877[ 1 ] = fresh_wire_874[ 1 ];
	assign fresh_wire_877[ 2 ] = fresh_wire_874[ 2 ];
	assign fresh_wire_877[ 3 ] = fresh_wire_874[ 3 ];
	assign fresh_wire_877[ 4 ] = fresh_wire_874[ 4 ];
	assign fresh_wire_877[ 5 ] = fresh_wire_874[ 5 ];
	assign fresh_wire_877[ 6 ] = fresh_wire_874[ 6 ];
	assign fresh_wire_877[ 7 ] = fresh_wire_874[ 7 ];
	assign fresh_wire_877[ 8 ] = fresh_wire_874[ 8 ];
	assign fresh_wire_877[ 9 ] = fresh_wire_874[ 9 ];
	assign fresh_wire_877[ 10 ] = fresh_wire_874[ 10 ];
	assign fresh_wire_877[ 11 ] = fresh_wire_874[ 11 ];
	assign fresh_wire_877[ 12 ] = fresh_wire_874[ 12 ];
	assign fresh_wire_877[ 13 ] = fresh_wire_874[ 13 ];
	assign fresh_wire_877[ 14 ] = fresh_wire_874[ 14 ];
	assign fresh_wire_877[ 15 ] = fresh_wire_874[ 15 ];
	assign fresh_wire_879[ 0 ] = fresh_wire_737[ 0 ];
	assign fresh_wire_880[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_881[ 0 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_883[ 0 ] = fresh_wire_826[ 0 ];
	assign fresh_wire_884[ 0 ] = fresh_wire_882[ 0 ];
	assign fresh_wire_885[ 0 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_887[ 0 ] = fresh_wire_819[ 0 ];
	assign fresh_wire_888[ 0 ] = fresh_wire_886[ 0 ];
	assign fresh_wire_889[ 0 ] = fresh_wire_758[ 0 ];
	assign fresh_wire_891[ 0 ] = fresh_wire_812[ 0 ];
	assign fresh_wire_892[ 0 ] = fresh_wire_890[ 0 ];
	assign fresh_wire_893[ 0 ] = fresh_wire_755[ 0 ];
	assign fresh_wire_895[ 0 ] = fresh_wire_798[ 0 ];
	assign fresh_wire_896[ 0 ] = fresh_wire_858[ 0 ];
	assign fresh_wire_896[ 1 ] = fresh_wire_858[ 1 ];
	assign fresh_wire_897[ 0 ] = fresh_wire_722[ 0 ];
	assign fresh_wire_897[ 1 ] = fresh_wire_722[ 1 ];
	assign fresh_wire_899[ 0 ] = fresh_wire_784[ 0 ];
	assign fresh_wire_900[ 0 ] = fresh_wire_898[ 0 ];
	assign fresh_wire_900[ 1 ] = fresh_wire_898[ 1 ];
	assign fresh_wire_901[ 0 ] = fresh_wire_858[ 0 ];
	assign fresh_wire_901[ 1 ] = fresh_wire_858[ 1 ];
	assign fresh_wire_903[ 0 ] = fresh_wire_777[ 0 ];
	assign fresh_wire_904[ 0 ] = fresh_wire_902[ 0 ];
	assign fresh_wire_904[ 1 ] = fresh_wire_902[ 1 ];
	assign fresh_wire_905[ 0 ] = fresh_wire_725[ 0 ];
	assign fresh_wire_905[ 1 ] = fresh_wire_725[ 1 ];
	assign fresh_wire_907[ 0 ] = fresh_wire_770[ 0 ];
	assign fresh_wire_908[ 0 ] = fresh_wire_906[ 0 ];
	assign fresh_wire_908[ 1 ] = fresh_wire_906[ 1 ];
	assign fresh_wire_909[ 0 ] = fresh_wire_722[ 0 ];
	assign fresh_wire_909[ 1 ] = fresh_wire_722[ 1 ];
	assign fresh_wire_911[ 0 ] = fresh_wire_763[ 0 ];
	assign fresh_wire_912[ 0 ] = fresh_wire_910[ 0 ];
	assign fresh_wire_912[ 1 ] = fresh_wire_910[ 1 ];
	assign fresh_wire_913[ 0 ] = fresh_wire_926[ 0 ];
	assign fresh_wire_913[ 1 ] = fresh_wire_926[ 1 ];
	assign fresh_wire_915[ 0 ] = fresh_wire_840[ 0 ];
	assign fresh_wire_916[ 0 ] = fresh_wire_862[ 0 ];
	assign fresh_wire_916[ 1 ] = fresh_wire_862[ 1 ];
	assign fresh_wire_916[ 2 ] = fresh_wire_862[ 2 ];
	assign fresh_wire_916[ 3 ] = fresh_wire_862[ 3 ];
	assign fresh_wire_916[ 4 ] = fresh_wire_862[ 4 ];
	assign fresh_wire_916[ 5 ] = fresh_wire_862[ 5 ];
	assign fresh_wire_916[ 6 ] = fresh_wire_862[ 6 ];
	assign fresh_wire_916[ 7 ] = fresh_wire_862[ 7 ];
	assign fresh_wire_916[ 8 ] = fresh_wire_862[ 8 ];
	assign fresh_wire_916[ 9 ] = fresh_wire_862[ 9 ];
	assign fresh_wire_916[ 10 ] = fresh_wire_862[ 10 ];
	assign fresh_wire_916[ 11 ] = fresh_wire_862[ 11 ];
	assign fresh_wire_916[ 12 ] = fresh_wire_862[ 12 ];
	assign fresh_wire_916[ 13 ] = fresh_wire_862[ 13 ];
	assign fresh_wire_916[ 14 ] = fresh_wire_862[ 14 ];
	assign fresh_wire_916[ 15 ] = fresh_wire_862[ 15 ];
	assign fresh_wire_916[ 16 ] = fresh_wire_862[ 16 ];
	assign fresh_wire_916[ 17 ] = fresh_wire_862[ 17 ];
	assign fresh_wire_916[ 18 ] = fresh_wire_862[ 18 ];
	assign fresh_wire_916[ 19 ] = fresh_wire_862[ 19 ];
	assign fresh_wire_916[ 20 ] = fresh_wire_862[ 20 ];
	assign fresh_wire_916[ 21 ] = fresh_wire_862[ 21 ];
	assign fresh_wire_916[ 22 ] = fresh_wire_862[ 22 ];
	assign fresh_wire_916[ 23 ] = fresh_wire_862[ 23 ];
	assign fresh_wire_916[ 24 ] = fresh_wire_862[ 24 ];
	assign fresh_wire_916[ 25 ] = fresh_wire_862[ 25 ];
	assign fresh_wire_916[ 26 ] = fresh_wire_862[ 26 ];
	assign fresh_wire_916[ 27 ] = fresh_wire_862[ 27 ];
	assign fresh_wire_916[ 28 ] = fresh_wire_862[ 28 ];
	assign fresh_wire_916[ 29 ] = fresh_wire_862[ 29 ];
	assign fresh_wire_916[ 30 ] = fresh_wire_862[ 30 ];
	assign fresh_wire_916[ 31 ] = fresh_wire_862[ 31 ];
	assign fresh_wire_916[ 32 ] = fresh_wire_862[ 32 ];
	assign fresh_wire_916[ 33 ] = fresh_wire_862[ 33 ];
	assign fresh_wire_916[ 34 ] = fresh_wire_862[ 34 ];
	assign fresh_wire_916[ 35 ] = fresh_wire_862[ 35 ];
	assign fresh_wire_916[ 36 ] = fresh_wire_862[ 36 ];
	assign fresh_wire_916[ 37 ] = fresh_wire_862[ 37 ];
	assign fresh_wire_916[ 38 ] = fresh_wire_862[ 38 ];
	assign fresh_wire_916[ 39 ] = fresh_wire_862[ 39 ];
	assign fresh_wire_916[ 40 ] = fresh_wire_862[ 40 ];
	assign fresh_wire_916[ 41 ] = fresh_wire_862[ 41 ];
	assign fresh_wire_916[ 42 ] = fresh_wire_862[ 42 ];
	assign fresh_wire_916[ 43 ] = fresh_wire_862[ 43 ];
	assign fresh_wire_916[ 44 ] = fresh_wire_862[ 44 ];
	assign fresh_wire_916[ 45 ] = fresh_wire_862[ 45 ];
	assign fresh_wire_916[ 46 ] = fresh_wire_862[ 46 ];
	assign fresh_wire_916[ 47 ] = fresh_wire_862[ 47 ];
	assign fresh_wire_917[ 0 ] = fresh_wire_600[ 0 ];
	assign fresh_wire_917[ 1 ] = fresh_wire_600[ 1 ];
	assign fresh_wire_917[ 2 ] = fresh_wire_600[ 2 ];
	assign fresh_wire_917[ 3 ] = fresh_wire_600[ 3 ];
	assign fresh_wire_917[ 4 ] = fresh_wire_600[ 4 ];
	assign fresh_wire_917[ 5 ] = fresh_wire_600[ 5 ];
	assign fresh_wire_917[ 6 ] = fresh_wire_600[ 6 ];
	assign fresh_wire_917[ 7 ] = fresh_wire_600[ 7 ];
	assign fresh_wire_917[ 8 ] = fresh_wire_600[ 8 ];
	assign fresh_wire_917[ 9 ] = fresh_wire_600[ 9 ];
	assign fresh_wire_917[ 10 ] = fresh_wire_600[ 10 ];
	assign fresh_wire_917[ 11 ] = fresh_wire_600[ 11 ];
	assign fresh_wire_917[ 12 ] = fresh_wire_600[ 12 ];
	assign fresh_wire_917[ 13 ] = fresh_wire_600[ 13 ];
	assign fresh_wire_917[ 14 ] = fresh_wire_600[ 14 ];
	assign fresh_wire_917[ 15 ] = fresh_wire_600[ 15 ];
	assign fresh_wire_917[ 16 ] = fresh_wire_862[ 0 ];
	assign fresh_wire_917[ 17 ] = fresh_wire_862[ 1 ];
	assign fresh_wire_917[ 18 ] = fresh_wire_862[ 2 ];
	assign fresh_wire_917[ 19 ] = fresh_wire_862[ 3 ];
	assign fresh_wire_917[ 20 ] = fresh_wire_862[ 4 ];
	assign fresh_wire_917[ 21 ] = fresh_wire_862[ 5 ];
	assign fresh_wire_917[ 22 ] = fresh_wire_862[ 6 ];
	assign fresh_wire_917[ 23 ] = fresh_wire_862[ 7 ];
	assign fresh_wire_917[ 24 ] = fresh_wire_862[ 8 ];
	assign fresh_wire_917[ 25 ] = fresh_wire_862[ 9 ];
	assign fresh_wire_917[ 26 ] = fresh_wire_862[ 10 ];
	assign fresh_wire_917[ 27 ] = fresh_wire_862[ 11 ];
	assign fresh_wire_917[ 28 ] = fresh_wire_862[ 12 ];
	assign fresh_wire_917[ 29 ] = fresh_wire_862[ 13 ];
	assign fresh_wire_917[ 30 ] = fresh_wire_862[ 14 ];
	assign fresh_wire_917[ 31 ] = fresh_wire_862[ 15 ];
	assign fresh_wire_917[ 32 ] = fresh_wire_862[ 16 ];
	assign fresh_wire_917[ 33 ] = fresh_wire_862[ 17 ];
	assign fresh_wire_917[ 34 ] = fresh_wire_862[ 18 ];
	assign fresh_wire_917[ 35 ] = fresh_wire_862[ 19 ];
	assign fresh_wire_917[ 36 ] = fresh_wire_862[ 20 ];
	assign fresh_wire_917[ 37 ] = fresh_wire_862[ 21 ];
	assign fresh_wire_917[ 38 ] = fresh_wire_862[ 22 ];
	assign fresh_wire_917[ 39 ] = fresh_wire_862[ 23 ];
	assign fresh_wire_917[ 40 ] = fresh_wire_862[ 24 ];
	assign fresh_wire_917[ 41 ] = fresh_wire_862[ 25 ];
	assign fresh_wire_917[ 42 ] = fresh_wire_862[ 26 ];
	assign fresh_wire_917[ 43 ] = fresh_wire_862[ 27 ];
	assign fresh_wire_917[ 44 ] = fresh_wire_862[ 28 ];
	assign fresh_wire_917[ 45 ] = fresh_wire_862[ 29 ];
	assign fresh_wire_917[ 46 ] = fresh_wire_862[ 30 ];
	assign fresh_wire_917[ 47 ] = fresh_wire_862[ 31 ];
	assign fresh_wire_919[ 0 ] = fresh_wire_728[ 0 ];
	assign fresh_wire_920[ 0 ] = fresh_wire_918[ 0 ];
	assign fresh_wire_920[ 1 ] = fresh_wire_918[ 1 ];
	assign fresh_wire_920[ 2 ] = fresh_wire_918[ 2 ];
	assign fresh_wire_920[ 3 ] = fresh_wire_918[ 3 ];
	assign fresh_wire_920[ 4 ] = fresh_wire_918[ 4 ];
	assign fresh_wire_920[ 5 ] = fresh_wire_918[ 5 ];
	assign fresh_wire_920[ 6 ] = fresh_wire_918[ 6 ];
	assign fresh_wire_920[ 7 ] = fresh_wire_918[ 7 ];
	assign fresh_wire_920[ 8 ] = fresh_wire_918[ 8 ];
	assign fresh_wire_920[ 9 ] = fresh_wire_918[ 9 ];
	assign fresh_wire_920[ 10 ] = fresh_wire_918[ 10 ];
	assign fresh_wire_920[ 11 ] = fresh_wire_918[ 11 ];
	assign fresh_wire_920[ 12 ] = fresh_wire_918[ 12 ];
	assign fresh_wire_920[ 13 ] = fresh_wire_918[ 13 ];
	assign fresh_wire_920[ 14 ] = fresh_wire_918[ 14 ];
	assign fresh_wire_920[ 15 ] = fresh_wire_918[ 15 ];
	assign fresh_wire_920[ 16 ] = fresh_wire_918[ 16 ];
	assign fresh_wire_920[ 17 ] = fresh_wire_918[ 17 ];
	assign fresh_wire_920[ 18 ] = fresh_wire_918[ 18 ];
	assign fresh_wire_920[ 19 ] = fresh_wire_918[ 19 ];
	assign fresh_wire_920[ 20 ] = fresh_wire_918[ 20 ];
	assign fresh_wire_920[ 21 ] = fresh_wire_918[ 21 ];
	assign fresh_wire_920[ 22 ] = fresh_wire_918[ 22 ];
	assign fresh_wire_920[ 23 ] = fresh_wire_918[ 23 ];
	assign fresh_wire_920[ 24 ] = fresh_wire_918[ 24 ];
	assign fresh_wire_920[ 25 ] = fresh_wire_918[ 25 ];
	assign fresh_wire_920[ 26 ] = fresh_wire_918[ 26 ];
	assign fresh_wire_920[ 27 ] = fresh_wire_918[ 27 ];
	assign fresh_wire_920[ 28 ] = fresh_wire_918[ 28 ];
	assign fresh_wire_920[ 29 ] = fresh_wire_918[ 29 ];
	assign fresh_wire_920[ 30 ] = fresh_wire_918[ 30 ];
	assign fresh_wire_920[ 31 ] = fresh_wire_918[ 31 ];
	assign fresh_wire_920[ 32 ] = fresh_wire_918[ 32 ];
	assign fresh_wire_920[ 33 ] = fresh_wire_918[ 33 ];
	assign fresh_wire_920[ 34 ] = fresh_wire_918[ 34 ];
	assign fresh_wire_920[ 35 ] = fresh_wire_918[ 35 ];
	assign fresh_wire_920[ 36 ] = fresh_wire_918[ 36 ];
	assign fresh_wire_920[ 37 ] = fresh_wire_918[ 37 ];
	assign fresh_wire_920[ 38 ] = fresh_wire_918[ 38 ];
	assign fresh_wire_920[ 39 ] = fresh_wire_918[ 39 ];
	assign fresh_wire_920[ 40 ] = fresh_wire_918[ 40 ];
	assign fresh_wire_920[ 41 ] = fresh_wire_918[ 41 ];
	assign fresh_wire_920[ 42 ] = fresh_wire_918[ 42 ];
	assign fresh_wire_920[ 43 ] = fresh_wire_918[ 43 ];
	assign fresh_wire_920[ 44 ] = fresh_wire_918[ 44 ];
	assign fresh_wire_920[ 45 ] = fresh_wire_918[ 45 ];
	assign fresh_wire_920[ 46 ] = fresh_wire_918[ 46 ];
	assign fresh_wire_920[ 47 ] = fresh_wire_918[ 47 ];
	assign fresh_wire_921[ 0 ] = fresh_wire_600[ 0 ];
	assign fresh_wire_921[ 1 ] = fresh_wire_600[ 1 ];
	assign fresh_wire_921[ 2 ] = fresh_wire_600[ 2 ];
	assign fresh_wire_921[ 3 ] = fresh_wire_600[ 3 ];
	assign fresh_wire_921[ 4 ] = fresh_wire_600[ 4 ];
	assign fresh_wire_921[ 5 ] = fresh_wire_600[ 5 ];
	assign fresh_wire_921[ 6 ] = fresh_wire_600[ 6 ];
	assign fresh_wire_921[ 7 ] = fresh_wire_600[ 7 ];
	assign fresh_wire_921[ 8 ] = fresh_wire_600[ 8 ];
	assign fresh_wire_921[ 9 ] = fresh_wire_600[ 9 ];
	assign fresh_wire_921[ 10 ] = fresh_wire_600[ 10 ];
	assign fresh_wire_921[ 11 ] = fresh_wire_600[ 11 ];
	assign fresh_wire_921[ 12 ] = fresh_wire_600[ 12 ];
	assign fresh_wire_921[ 13 ] = fresh_wire_600[ 13 ];
	assign fresh_wire_921[ 14 ] = fresh_wire_600[ 14 ];
	assign fresh_wire_921[ 15 ] = fresh_wire_600[ 15 ];
	assign fresh_wire_921[ 16 ] = fresh_wire_600[ 16 ];
	assign fresh_wire_921[ 17 ] = fresh_wire_600[ 17 ];
	assign fresh_wire_921[ 18 ] = fresh_wire_600[ 18 ];
	assign fresh_wire_921[ 19 ] = fresh_wire_600[ 19 ];
	assign fresh_wire_921[ 20 ] = fresh_wire_600[ 20 ];
	assign fresh_wire_921[ 21 ] = fresh_wire_600[ 21 ];
	assign fresh_wire_921[ 22 ] = fresh_wire_600[ 22 ];
	assign fresh_wire_921[ 23 ] = fresh_wire_600[ 23 ];
	assign fresh_wire_921[ 24 ] = fresh_wire_600[ 24 ];
	assign fresh_wire_921[ 25 ] = fresh_wire_600[ 25 ];
	assign fresh_wire_921[ 26 ] = fresh_wire_600[ 26 ];
	assign fresh_wire_921[ 27 ] = fresh_wire_600[ 27 ];
	assign fresh_wire_921[ 28 ] = fresh_wire_600[ 28 ];
	assign fresh_wire_921[ 29 ] = fresh_wire_600[ 29 ];
	assign fresh_wire_921[ 30 ] = fresh_wire_600[ 30 ];
	assign fresh_wire_921[ 31 ] = fresh_wire_600[ 31 ];
	assign fresh_wire_921[ 32 ] = fresh_wire_862[ 0 ];
	assign fresh_wire_921[ 33 ] = fresh_wire_862[ 1 ];
	assign fresh_wire_921[ 34 ] = fresh_wire_862[ 2 ];
	assign fresh_wire_921[ 35 ] = fresh_wire_862[ 3 ];
	assign fresh_wire_921[ 36 ] = fresh_wire_862[ 4 ];
	assign fresh_wire_921[ 37 ] = fresh_wire_862[ 5 ];
	assign fresh_wire_921[ 38 ] = fresh_wire_862[ 6 ];
	assign fresh_wire_921[ 39 ] = fresh_wire_862[ 7 ];
	assign fresh_wire_921[ 40 ] = fresh_wire_862[ 8 ];
	assign fresh_wire_921[ 41 ] = fresh_wire_862[ 9 ];
	assign fresh_wire_921[ 42 ] = fresh_wire_862[ 10 ];
	assign fresh_wire_921[ 43 ] = fresh_wire_862[ 11 ];
	assign fresh_wire_921[ 44 ] = fresh_wire_862[ 12 ];
	assign fresh_wire_921[ 45 ] = fresh_wire_862[ 13 ];
	assign fresh_wire_921[ 46 ] = fresh_wire_862[ 14 ];
	assign fresh_wire_921[ 47 ] = fresh_wire_862[ 15 ];
	assign fresh_wire_923[ 0 ] = fresh_wire_734[ 0 ];
	assign fresh_wire_924[ 0 ] = fresh_wire_858[ 0 ];
	assign fresh_wire_924[ 1 ] = fresh_wire_858[ 1 ];
	assign fresh_wire_925[ 0 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_925[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_928[ 0 ] = fresh_wire_157[ 0 ];
	assign fresh_wire_930[ 0 ] = fresh_wire_426[ 0 ];
	assign fresh_wire_932[ 0 ] = fresh_wire_929[ 0 ];
	assign fresh_wire_933[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_935[ 0 ] = fresh_wire_931[ 0 ];
	assign fresh_wire_936[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_938[ 0 ] = fresh_wire_943[ 0 ];
	assign fresh_wire_938[ 1 ] = fresh_wire_943[ 1 ];
	assign fresh_wire_938[ 2 ] = fresh_wire_943[ 2 ];
	assign fresh_wire_938[ 3 ] = fresh_wire_943[ 3 ];
	assign fresh_wire_938[ 4 ] = fresh_wire_943[ 4 ];
	assign fresh_wire_938[ 5 ] = fresh_wire_943[ 5 ];
	assign fresh_wire_938[ 6 ] = fresh_wire_943[ 6 ];
	assign fresh_wire_938[ 7 ] = fresh_wire_943[ 7 ];
	assign fresh_wire_938[ 8 ] = fresh_wire_943[ 8 ];
	assign fresh_wire_938[ 9 ] = fresh_wire_943[ 9 ];
	assign fresh_wire_938[ 10 ] = fresh_wire_943[ 10 ];
	assign fresh_wire_938[ 11 ] = fresh_wire_943[ 11 ];
	assign fresh_wire_938[ 12 ] = fresh_wire_943[ 12 ];
	assign fresh_wire_938[ 13 ] = fresh_wire_943[ 13 ];
	assign fresh_wire_938[ 14 ] = fresh_wire_943[ 14 ];
	assign fresh_wire_938[ 15 ] = fresh_wire_943[ 15 ];
	assign fresh_wire_940[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_941[ 0 ] = fresh_wire_939[ 0 ];
	assign fresh_wire_941[ 1 ] = fresh_wire_939[ 1 ];
	assign fresh_wire_941[ 2 ] = fresh_wire_939[ 2 ];
	assign fresh_wire_941[ 3 ] = fresh_wire_939[ 3 ];
	assign fresh_wire_941[ 4 ] = fresh_wire_939[ 4 ];
	assign fresh_wire_941[ 5 ] = fresh_wire_939[ 5 ];
	assign fresh_wire_941[ 6 ] = fresh_wire_939[ 6 ];
	assign fresh_wire_941[ 7 ] = fresh_wire_939[ 7 ];
	assign fresh_wire_941[ 8 ] = fresh_wire_939[ 8 ];
	assign fresh_wire_941[ 9 ] = fresh_wire_939[ 9 ];
	assign fresh_wire_941[ 10 ] = fresh_wire_939[ 10 ];
	assign fresh_wire_941[ 11 ] = fresh_wire_939[ 11 ];
	assign fresh_wire_941[ 12 ] = fresh_wire_939[ 12 ];
	assign fresh_wire_941[ 13 ] = fresh_wire_939[ 13 ];
	assign fresh_wire_941[ 14 ] = fresh_wire_939[ 14 ];
	assign fresh_wire_941[ 15 ] = fresh_wire_939[ 15 ];
	assign fresh_wire_942[ 0 ] = fresh_wire_1022[ 0 ];
	assign fresh_wire_942[ 1 ] = fresh_wire_1022[ 1 ];
	assign fresh_wire_942[ 2 ] = fresh_wire_1022[ 2 ];
	assign fresh_wire_942[ 3 ] = fresh_wire_1022[ 3 ];
	assign fresh_wire_942[ 4 ] = fresh_wire_1022[ 4 ];
	assign fresh_wire_942[ 5 ] = fresh_wire_1022[ 5 ];
	assign fresh_wire_942[ 6 ] = fresh_wire_1022[ 6 ];
	assign fresh_wire_942[ 7 ] = fresh_wire_1022[ 7 ];
	assign fresh_wire_942[ 8 ] = fresh_wire_1022[ 8 ];
	assign fresh_wire_942[ 9 ] = fresh_wire_1022[ 9 ];
	assign fresh_wire_942[ 10 ] = fresh_wire_1022[ 10 ];
	assign fresh_wire_942[ 11 ] = fresh_wire_1022[ 11 ];
	assign fresh_wire_942[ 12 ] = fresh_wire_1022[ 12 ];
	assign fresh_wire_942[ 13 ] = fresh_wire_1022[ 13 ];
	assign fresh_wire_942[ 14 ] = fresh_wire_1022[ 14 ];
	assign fresh_wire_942[ 15 ] = fresh_wire_1022[ 15 ];
	assign fresh_wire_944[ 0 ] = fresh_wire_934[ 0 ];
	assign fresh_wire_945[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_945[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_945[ 2 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_945[ 3 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_945[ 4 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_945[ 5 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_945[ 6 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_945[ 7 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_945[ 8 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_945[ 9 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_945[ 10 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_945[ 11 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_945[ 12 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_945[ 13 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_945[ 14 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_945[ 15 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_946[ 0 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 1 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 2 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 3 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 4 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 5 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 6 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 7 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 8 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 9 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 10 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 11 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 12 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 13 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 14 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 15 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_948[ 0 ] = fresh_wire_937[ 0 ];
	assign fresh_wire_950[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_950[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_950[ 2 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_950[ 3 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_950[ 4 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_950[ 5 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_950[ 6 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_950[ 7 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_950[ 8 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_950[ 9 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_950[ 10 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_950[ 11 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_950[ 12 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_950[ 13 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_950[ 14 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_950[ 15 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_951[ 0 ] = fresh_wire_947[ 0 ];
	assign fresh_wire_951[ 1 ] = fresh_wire_947[ 1 ];
	assign fresh_wire_951[ 2 ] = fresh_wire_947[ 2 ];
	assign fresh_wire_951[ 3 ] = fresh_wire_947[ 3 ];
	assign fresh_wire_951[ 4 ] = fresh_wire_947[ 4 ];
	assign fresh_wire_951[ 5 ] = fresh_wire_947[ 5 ];
	assign fresh_wire_951[ 6 ] = fresh_wire_947[ 6 ];
	assign fresh_wire_951[ 7 ] = fresh_wire_947[ 7 ];
	assign fresh_wire_951[ 8 ] = fresh_wire_947[ 8 ];
	assign fresh_wire_951[ 9 ] = fresh_wire_947[ 9 ];
	assign fresh_wire_951[ 10 ] = fresh_wire_947[ 10 ];
	assign fresh_wire_951[ 11 ] = fresh_wire_947[ 11 ];
	assign fresh_wire_951[ 12 ] = fresh_wire_947[ 12 ];
	assign fresh_wire_951[ 13 ] = fresh_wire_947[ 13 ];
	assign fresh_wire_951[ 14 ] = fresh_wire_947[ 14 ];
	assign fresh_wire_951[ 15 ] = fresh_wire_947[ 15 ];
	assign fresh_wire_953[ 0 ] = fresh_wire_934[ 0 ];
	assign fresh_wire_954[ 0 ] = fresh_wire_958[ 0 ];
	assign fresh_wire_954[ 1 ] = fresh_wire_965[ 0 ];
	assign fresh_wire_954[ 2 ] = fresh_wire_966[ 0 ];
	assign fresh_wire_954[ 3 ] = fresh_wire_967[ 0 ];
	assign fresh_wire_954[ 4 ] = fresh_wire_968[ 0 ];
	assign fresh_wire_954[ 5 ] = fresh_wire_969[ 0 ];
	assign fresh_wire_954[ 6 ] = fresh_wire_970[ 0 ];
	assign fresh_wire_954[ 7 ] = fresh_wire_971[ 0 ];
	assign fresh_wire_954[ 8 ] = fresh_wire_972[ 0 ];
	assign fresh_wire_954[ 9 ] = fresh_wire_973[ 0 ];
	assign fresh_wire_954[ 10 ] = fresh_wire_959[ 0 ];
	assign fresh_wire_954[ 11 ] = fresh_wire_960[ 0 ];
	assign fresh_wire_954[ 12 ] = fresh_wire_961[ 0 ];
	assign fresh_wire_954[ 13 ] = fresh_wire_962[ 0 ];
	assign fresh_wire_954[ 14 ] = fresh_wire_963[ 0 ];
	assign fresh_wire_954[ 15 ] = fresh_wire_964[ 0 ];
	assign fresh_wire_955[ 0 ] = fresh_wire_714[ 0 ];
	assign fresh_wire_955[ 1 ] = fresh_wire_714[ 1 ];
	assign fresh_wire_955[ 2 ] = fresh_wire_714[ 2 ];
	assign fresh_wire_955[ 3 ] = fresh_wire_714[ 3 ];
	assign fresh_wire_955[ 4 ] = fresh_wire_714[ 4 ];
	assign fresh_wire_955[ 5 ] = fresh_wire_714[ 5 ];
	assign fresh_wire_955[ 6 ] = fresh_wire_714[ 6 ];
	assign fresh_wire_955[ 7 ] = fresh_wire_714[ 7 ];
	assign fresh_wire_955[ 8 ] = fresh_wire_714[ 8 ];
	assign fresh_wire_955[ 9 ] = fresh_wire_714[ 9 ];
	assign fresh_wire_955[ 10 ] = fresh_wire_714[ 10 ];
	assign fresh_wire_955[ 11 ] = fresh_wire_714[ 11 ];
	assign fresh_wire_955[ 12 ] = fresh_wire_714[ 12 ];
	assign fresh_wire_955[ 13 ] = fresh_wire_714[ 13 ];
	assign fresh_wire_955[ 14 ] = fresh_wire_714[ 14 ];
	assign fresh_wire_955[ 15 ] = fresh_wire_714[ 15 ];
	assign fresh_wire_957[ 0 ] = fresh_wire_937[ 0 ];
	assign fresh_wire_974[ 0 ] = fresh_wire_978[ 0 ];
	assign fresh_wire_974[ 1 ] = fresh_wire_985[ 0 ];
	assign fresh_wire_974[ 2 ] = fresh_wire_986[ 0 ];
	assign fresh_wire_974[ 3 ] = fresh_wire_987[ 0 ];
	assign fresh_wire_974[ 4 ] = fresh_wire_988[ 0 ];
	assign fresh_wire_974[ 5 ] = fresh_wire_989[ 0 ];
	assign fresh_wire_974[ 6 ] = fresh_wire_990[ 0 ];
	assign fresh_wire_974[ 7 ] = fresh_wire_991[ 0 ];
	assign fresh_wire_974[ 8 ] = fresh_wire_992[ 0 ];
	assign fresh_wire_974[ 9 ] = fresh_wire_993[ 0 ];
	assign fresh_wire_974[ 10 ] = fresh_wire_979[ 0 ];
	assign fresh_wire_974[ 11 ] = fresh_wire_980[ 0 ];
	assign fresh_wire_974[ 12 ] = fresh_wire_981[ 0 ];
	assign fresh_wire_974[ 13 ] = fresh_wire_982[ 0 ];
	assign fresh_wire_974[ 14 ] = fresh_wire_983[ 0 ];
	assign fresh_wire_974[ 15 ] = fresh_wire_984[ 0 ];
	assign fresh_wire_975[ 0 ] = fresh_wire_956[ 0 ];
	assign fresh_wire_975[ 1 ] = fresh_wire_956[ 1 ];
	assign fresh_wire_975[ 2 ] = fresh_wire_956[ 2 ];
	assign fresh_wire_975[ 3 ] = fresh_wire_956[ 3 ];
	assign fresh_wire_975[ 4 ] = fresh_wire_956[ 4 ];
	assign fresh_wire_975[ 5 ] = fresh_wire_956[ 5 ];
	assign fresh_wire_975[ 6 ] = fresh_wire_956[ 6 ];
	assign fresh_wire_975[ 7 ] = fresh_wire_956[ 7 ];
	assign fresh_wire_975[ 8 ] = fresh_wire_956[ 8 ];
	assign fresh_wire_975[ 9 ] = fresh_wire_956[ 9 ];
	assign fresh_wire_975[ 10 ] = fresh_wire_956[ 10 ];
	assign fresh_wire_975[ 11 ] = fresh_wire_956[ 11 ];
	assign fresh_wire_975[ 12 ] = fresh_wire_956[ 12 ];
	assign fresh_wire_975[ 13 ] = fresh_wire_956[ 13 ];
	assign fresh_wire_975[ 14 ] = fresh_wire_956[ 14 ];
	assign fresh_wire_975[ 15 ] = fresh_wire_956[ 15 ];
	assign fresh_wire_977[ 0 ] = fresh_wire_934[ 0 ];
	assign fresh_wire_994[ 0 ] = fresh_wire_998[ 0 ];
	assign fresh_wire_994[ 1 ] = fresh_wire_999[ 0 ];
	assign fresh_wire_994[ 2 ] = fresh_wire_1000[ 0 ];
	assign fresh_wire_994[ 3 ] = fresh_wire_1001[ 0 ];
	assign fresh_wire_994[ 4 ] = fresh_wire_1002[ 0 ];
	assign fresh_wire_994[ 5 ] = fresh_wire_1003[ 0 ];
	assign fresh_wire_994[ 6 ] = fresh_wire_1004[ 0 ];
	assign fresh_wire_994[ 7 ] = fresh_wire_1005[ 0 ];
	assign fresh_wire_994[ 8 ] = fresh_wire_1006[ 0 ];
	assign fresh_wire_995[ 0 ] = fresh_wire_435[ 0 ];
	assign fresh_wire_995[ 1 ] = fresh_wire_435[ 1 ];
	assign fresh_wire_995[ 2 ] = fresh_wire_435[ 2 ];
	assign fresh_wire_995[ 3 ] = fresh_wire_435[ 3 ];
	assign fresh_wire_995[ 4 ] = fresh_wire_435[ 4 ];
	assign fresh_wire_995[ 5 ] = fresh_wire_435[ 5 ];
	assign fresh_wire_995[ 6 ] = fresh_wire_435[ 6 ];
	assign fresh_wire_995[ 7 ] = fresh_wire_435[ 7 ];
	assign fresh_wire_995[ 8 ] = fresh_wire_435[ 8 ];
	assign fresh_wire_997[ 0 ] = fresh_wire_937[ 0 ];
	assign fresh_wire_1007[ 0 ] = fresh_wire_1011[ 0 ];
	assign fresh_wire_1007[ 1 ] = fresh_wire_1012[ 0 ];
	assign fresh_wire_1007[ 2 ] = fresh_wire_1013[ 0 ];
	assign fresh_wire_1007[ 3 ] = fresh_wire_1014[ 0 ];
	assign fresh_wire_1007[ 4 ] = fresh_wire_1015[ 0 ];
	assign fresh_wire_1007[ 5 ] = fresh_wire_1016[ 0 ];
	assign fresh_wire_1007[ 6 ] = fresh_wire_1017[ 0 ];
	assign fresh_wire_1007[ 7 ] = fresh_wire_1018[ 0 ];
	assign fresh_wire_1007[ 8 ] = fresh_wire_1019[ 0 ];
	assign fresh_wire_1008[ 0 ] = fresh_wire_996[ 0 ];
	assign fresh_wire_1008[ 1 ] = fresh_wire_996[ 1 ];
	assign fresh_wire_1008[ 2 ] = fresh_wire_996[ 2 ];
	assign fresh_wire_1008[ 3 ] = fresh_wire_996[ 3 ];
	assign fresh_wire_1008[ 4 ] = fresh_wire_996[ 4 ];
	assign fresh_wire_1008[ 5 ] = fresh_wire_996[ 5 ];
	assign fresh_wire_1008[ 6 ] = fresh_wire_996[ 6 ];
	assign fresh_wire_1008[ 7 ] = fresh_wire_996[ 7 ];
	assign fresh_wire_1008[ 8 ] = fresh_wire_996[ 8 ];
	assign fresh_wire_1010[ 0 ] = fresh_wire_934[ 0 ];
	assign fresh_wire_1020[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1021[ 0 ] = fresh_wire_435[ 0 ];
	assign fresh_wire_1021[ 1 ] = fresh_wire_435[ 1 ];
	assign fresh_wire_1021[ 2 ] = fresh_wire_435[ 2 ];
	assign fresh_wire_1021[ 3 ] = fresh_wire_435[ 3 ];
	assign fresh_wire_1021[ 4 ] = fresh_wire_435[ 4 ];
	assign fresh_wire_1021[ 5 ] = fresh_wire_435[ 5 ];
	assign fresh_wire_1021[ 6 ] = fresh_wire_435[ 6 ];
	assign fresh_wire_1021[ 7 ] = fresh_wire_435[ 7 ];
	assign fresh_wire_1021[ 8 ] = fresh_wire_435[ 8 ];
	assign fresh_wire_1023[ 0 ] = fresh_wire_1009[ 0 ];
	assign fresh_wire_1023[ 1 ] = fresh_wire_1009[ 1 ];
	assign fresh_wire_1023[ 2 ] = fresh_wire_1009[ 2 ];
	assign fresh_wire_1023[ 3 ] = fresh_wire_1009[ 3 ];
	assign fresh_wire_1023[ 4 ] = fresh_wire_1009[ 4 ];
	assign fresh_wire_1023[ 5 ] = fresh_wire_1009[ 5 ];
	assign fresh_wire_1023[ 6 ] = fresh_wire_1009[ 6 ];
	assign fresh_wire_1023[ 7 ] = fresh_wire_1009[ 7 ];
	assign fresh_wire_1023[ 8 ] = fresh_wire_1009[ 8 ];
	assign fresh_wire_1024[ 0 ] = fresh_wire_976[ 0 ];
	assign fresh_wire_1024[ 1 ] = fresh_wire_976[ 1 ];
	assign fresh_wire_1024[ 2 ] = fresh_wire_976[ 2 ];
	assign fresh_wire_1024[ 3 ] = fresh_wire_976[ 3 ];
	assign fresh_wire_1024[ 4 ] = fresh_wire_976[ 4 ];
	assign fresh_wire_1024[ 5 ] = fresh_wire_976[ 5 ];
	assign fresh_wire_1024[ 6 ] = fresh_wire_976[ 6 ];
	assign fresh_wire_1024[ 7 ] = fresh_wire_976[ 7 ];
	assign fresh_wire_1024[ 8 ] = fresh_wire_976[ 8 ];
	assign fresh_wire_1024[ 9 ] = fresh_wire_976[ 9 ];
	assign fresh_wire_1024[ 10 ] = fresh_wire_976[ 10 ];
	assign fresh_wire_1024[ 11 ] = fresh_wire_976[ 11 ];
	assign fresh_wire_1024[ 12 ] = fresh_wire_976[ 12 ];
	assign fresh_wire_1024[ 13 ] = fresh_wire_976[ 13 ];
	assign fresh_wire_1024[ 14 ] = fresh_wire_976[ 14 ];
	assign fresh_wire_1024[ 15 ] = fresh_wire_976[ 15 ];
	assign fresh_wire_1025[ 0 ] = fresh_wire_952[ 0 ];
	assign fresh_wire_1026[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_1028[ 0 ] = fresh_wire_426[ 0 ];
	assign fresh_wire_1030[ 0 ] = fresh_wire_1027[ 0 ];
	assign fresh_wire_1031[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1033[ 0 ] = fresh_wire_1029[ 0 ];
	assign fresh_wire_1034[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1036[ 0 ] = fresh_wire_1041[ 0 ];
	assign fresh_wire_1036[ 1 ] = fresh_wire_1041[ 1 ];
	assign fresh_wire_1036[ 2 ] = fresh_wire_1041[ 2 ];
	assign fresh_wire_1036[ 3 ] = fresh_wire_1041[ 3 ];
	assign fresh_wire_1036[ 4 ] = fresh_wire_1041[ 4 ];
	assign fresh_wire_1036[ 5 ] = fresh_wire_1041[ 5 ];
	assign fresh_wire_1036[ 6 ] = fresh_wire_1041[ 6 ];
	assign fresh_wire_1036[ 7 ] = fresh_wire_1041[ 7 ];
	assign fresh_wire_1036[ 8 ] = fresh_wire_1041[ 8 ];
	assign fresh_wire_1036[ 9 ] = fresh_wire_1041[ 9 ];
	assign fresh_wire_1036[ 10 ] = fresh_wire_1041[ 10 ];
	assign fresh_wire_1036[ 11 ] = fresh_wire_1041[ 11 ];
	assign fresh_wire_1036[ 12 ] = fresh_wire_1041[ 12 ];
	assign fresh_wire_1036[ 13 ] = fresh_wire_1041[ 13 ];
	assign fresh_wire_1036[ 14 ] = fresh_wire_1041[ 14 ];
	assign fresh_wire_1036[ 15 ] = fresh_wire_1041[ 15 ];
	assign fresh_wire_1038[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1039[ 0 ] = fresh_wire_1037[ 0 ];
	assign fresh_wire_1039[ 1 ] = fresh_wire_1037[ 1 ];
	assign fresh_wire_1039[ 2 ] = fresh_wire_1037[ 2 ];
	assign fresh_wire_1039[ 3 ] = fresh_wire_1037[ 3 ];
	assign fresh_wire_1039[ 4 ] = fresh_wire_1037[ 4 ];
	assign fresh_wire_1039[ 5 ] = fresh_wire_1037[ 5 ];
	assign fresh_wire_1039[ 6 ] = fresh_wire_1037[ 6 ];
	assign fresh_wire_1039[ 7 ] = fresh_wire_1037[ 7 ];
	assign fresh_wire_1039[ 8 ] = fresh_wire_1037[ 8 ];
	assign fresh_wire_1039[ 9 ] = fresh_wire_1037[ 9 ];
	assign fresh_wire_1039[ 10 ] = fresh_wire_1037[ 10 ];
	assign fresh_wire_1039[ 11 ] = fresh_wire_1037[ 11 ];
	assign fresh_wire_1039[ 12 ] = fresh_wire_1037[ 12 ];
	assign fresh_wire_1039[ 13 ] = fresh_wire_1037[ 13 ];
	assign fresh_wire_1039[ 14 ] = fresh_wire_1037[ 14 ];
	assign fresh_wire_1039[ 15 ] = fresh_wire_1037[ 15 ];
	assign fresh_wire_1040[ 0 ] = fresh_wire_1120[ 0 ];
	assign fresh_wire_1040[ 1 ] = fresh_wire_1120[ 1 ];
	assign fresh_wire_1040[ 2 ] = fresh_wire_1120[ 2 ];
	assign fresh_wire_1040[ 3 ] = fresh_wire_1120[ 3 ];
	assign fresh_wire_1040[ 4 ] = fresh_wire_1120[ 4 ];
	assign fresh_wire_1040[ 5 ] = fresh_wire_1120[ 5 ];
	assign fresh_wire_1040[ 6 ] = fresh_wire_1120[ 6 ];
	assign fresh_wire_1040[ 7 ] = fresh_wire_1120[ 7 ];
	assign fresh_wire_1040[ 8 ] = fresh_wire_1120[ 8 ];
	assign fresh_wire_1040[ 9 ] = fresh_wire_1120[ 9 ];
	assign fresh_wire_1040[ 10 ] = fresh_wire_1120[ 10 ];
	assign fresh_wire_1040[ 11 ] = fresh_wire_1120[ 11 ];
	assign fresh_wire_1040[ 12 ] = fresh_wire_1120[ 12 ];
	assign fresh_wire_1040[ 13 ] = fresh_wire_1120[ 13 ];
	assign fresh_wire_1040[ 14 ] = fresh_wire_1120[ 14 ];
	assign fresh_wire_1040[ 15 ] = fresh_wire_1120[ 15 ];
	assign fresh_wire_1042[ 0 ] = fresh_wire_1032[ 0 ];
	assign fresh_wire_1043[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1043[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1043[ 2 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1043[ 3 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1043[ 4 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1043[ 5 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1043[ 6 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1043[ 7 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1043[ 8 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1043[ 9 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1043[ 10 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1043[ 11 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1043[ 12 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1043[ 13 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1043[ 14 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1043[ 15 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1044[ 0 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 1 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 2 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 3 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 4 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 5 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 6 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 7 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 8 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 9 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 10 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 11 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 12 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 13 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 14 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 15 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1046[ 0 ] = fresh_wire_1035[ 0 ];
	assign fresh_wire_1048[ 0 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1048[ 1 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1048[ 2 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1048[ 3 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1048[ 4 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1048[ 5 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1048[ 6 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1048[ 7 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1048[ 8 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1048[ 9 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1048[ 10 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1048[ 11 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1048[ 12 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1048[ 13 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1048[ 14 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1048[ 15 ] = fresh_wire_1152[ 0 ];
	assign fresh_wire_1049[ 0 ] = fresh_wire_1045[ 0 ];
	assign fresh_wire_1049[ 1 ] = fresh_wire_1045[ 1 ];
	assign fresh_wire_1049[ 2 ] = fresh_wire_1045[ 2 ];
	assign fresh_wire_1049[ 3 ] = fresh_wire_1045[ 3 ];
	assign fresh_wire_1049[ 4 ] = fresh_wire_1045[ 4 ];
	assign fresh_wire_1049[ 5 ] = fresh_wire_1045[ 5 ];
	assign fresh_wire_1049[ 6 ] = fresh_wire_1045[ 6 ];
	assign fresh_wire_1049[ 7 ] = fresh_wire_1045[ 7 ];
	assign fresh_wire_1049[ 8 ] = fresh_wire_1045[ 8 ];
	assign fresh_wire_1049[ 9 ] = fresh_wire_1045[ 9 ];
	assign fresh_wire_1049[ 10 ] = fresh_wire_1045[ 10 ];
	assign fresh_wire_1049[ 11 ] = fresh_wire_1045[ 11 ];
	assign fresh_wire_1049[ 12 ] = fresh_wire_1045[ 12 ];
	assign fresh_wire_1049[ 13 ] = fresh_wire_1045[ 13 ];
	assign fresh_wire_1049[ 14 ] = fresh_wire_1045[ 14 ];
	assign fresh_wire_1049[ 15 ] = fresh_wire_1045[ 15 ];
	assign fresh_wire_1051[ 0 ] = fresh_wire_1032[ 0 ];
	assign fresh_wire_1052[ 0 ] = fresh_wire_1056[ 0 ];
	assign fresh_wire_1052[ 1 ] = fresh_wire_1063[ 0 ];
	assign fresh_wire_1052[ 2 ] = fresh_wire_1064[ 0 ];
	assign fresh_wire_1052[ 3 ] = fresh_wire_1065[ 0 ];
	assign fresh_wire_1052[ 4 ] = fresh_wire_1066[ 0 ];
	assign fresh_wire_1052[ 5 ] = fresh_wire_1067[ 0 ];
	assign fresh_wire_1052[ 6 ] = fresh_wire_1068[ 0 ];
	assign fresh_wire_1052[ 7 ] = fresh_wire_1069[ 0 ];
	assign fresh_wire_1052[ 8 ] = fresh_wire_1070[ 0 ];
	assign fresh_wire_1052[ 9 ] = fresh_wire_1071[ 0 ];
	assign fresh_wire_1052[ 10 ] = fresh_wire_1057[ 0 ];
	assign fresh_wire_1052[ 11 ] = fresh_wire_1058[ 0 ];
	assign fresh_wire_1052[ 12 ] = fresh_wire_1059[ 0 ];
	assign fresh_wire_1052[ 13 ] = fresh_wire_1060[ 0 ];
	assign fresh_wire_1052[ 14 ] = fresh_wire_1061[ 0 ];
	assign fresh_wire_1052[ 15 ] = fresh_wire_1062[ 0 ];
	assign fresh_wire_1053[ 0 ] = fresh_wire_714[ 16 ];
	assign fresh_wire_1053[ 1 ] = fresh_wire_714[ 17 ];
	assign fresh_wire_1053[ 2 ] = fresh_wire_714[ 18 ];
	assign fresh_wire_1053[ 3 ] = fresh_wire_714[ 19 ];
	assign fresh_wire_1053[ 4 ] = fresh_wire_714[ 20 ];
	assign fresh_wire_1053[ 5 ] = fresh_wire_714[ 21 ];
	assign fresh_wire_1053[ 6 ] = fresh_wire_714[ 22 ];
	assign fresh_wire_1053[ 7 ] = fresh_wire_714[ 23 ];
	assign fresh_wire_1053[ 8 ] = fresh_wire_714[ 24 ];
	assign fresh_wire_1053[ 9 ] = fresh_wire_714[ 25 ];
	assign fresh_wire_1053[ 10 ] = fresh_wire_714[ 26 ];
	assign fresh_wire_1053[ 11 ] = fresh_wire_714[ 27 ];
	assign fresh_wire_1053[ 12 ] = fresh_wire_714[ 28 ];
	assign fresh_wire_1053[ 13 ] = fresh_wire_714[ 29 ];
	assign fresh_wire_1053[ 14 ] = fresh_wire_714[ 30 ];
	assign fresh_wire_1053[ 15 ] = fresh_wire_714[ 31 ];
	assign fresh_wire_1055[ 0 ] = fresh_wire_1035[ 0 ];
	assign fresh_wire_1072[ 0 ] = fresh_wire_1076[ 0 ];
	assign fresh_wire_1072[ 1 ] = fresh_wire_1083[ 0 ];
	assign fresh_wire_1072[ 2 ] = fresh_wire_1084[ 0 ];
	assign fresh_wire_1072[ 3 ] = fresh_wire_1085[ 0 ];
	assign fresh_wire_1072[ 4 ] = fresh_wire_1086[ 0 ];
	assign fresh_wire_1072[ 5 ] = fresh_wire_1087[ 0 ];
	assign fresh_wire_1072[ 6 ] = fresh_wire_1088[ 0 ];
	assign fresh_wire_1072[ 7 ] = fresh_wire_1089[ 0 ];
	assign fresh_wire_1072[ 8 ] = fresh_wire_1090[ 0 ];
	assign fresh_wire_1072[ 9 ] = fresh_wire_1091[ 0 ];
	assign fresh_wire_1072[ 10 ] = fresh_wire_1077[ 0 ];
	assign fresh_wire_1072[ 11 ] = fresh_wire_1078[ 0 ];
	assign fresh_wire_1072[ 12 ] = fresh_wire_1079[ 0 ];
	assign fresh_wire_1072[ 13 ] = fresh_wire_1080[ 0 ];
	assign fresh_wire_1072[ 14 ] = fresh_wire_1081[ 0 ];
	assign fresh_wire_1072[ 15 ] = fresh_wire_1082[ 0 ];
	assign fresh_wire_1073[ 0 ] = fresh_wire_1054[ 0 ];
	assign fresh_wire_1073[ 1 ] = fresh_wire_1054[ 1 ];
	assign fresh_wire_1073[ 2 ] = fresh_wire_1054[ 2 ];
	assign fresh_wire_1073[ 3 ] = fresh_wire_1054[ 3 ];
	assign fresh_wire_1073[ 4 ] = fresh_wire_1054[ 4 ];
	assign fresh_wire_1073[ 5 ] = fresh_wire_1054[ 5 ];
	assign fresh_wire_1073[ 6 ] = fresh_wire_1054[ 6 ];
	assign fresh_wire_1073[ 7 ] = fresh_wire_1054[ 7 ];
	assign fresh_wire_1073[ 8 ] = fresh_wire_1054[ 8 ];
	assign fresh_wire_1073[ 9 ] = fresh_wire_1054[ 9 ];
	assign fresh_wire_1073[ 10 ] = fresh_wire_1054[ 10 ];
	assign fresh_wire_1073[ 11 ] = fresh_wire_1054[ 11 ];
	assign fresh_wire_1073[ 12 ] = fresh_wire_1054[ 12 ];
	assign fresh_wire_1073[ 13 ] = fresh_wire_1054[ 13 ];
	assign fresh_wire_1073[ 14 ] = fresh_wire_1054[ 14 ];
	assign fresh_wire_1073[ 15 ] = fresh_wire_1054[ 15 ];
	assign fresh_wire_1075[ 0 ] = fresh_wire_1032[ 0 ];
	assign fresh_wire_1092[ 0 ] = fresh_wire_1096[ 0 ];
	assign fresh_wire_1092[ 1 ] = fresh_wire_1097[ 0 ];
	assign fresh_wire_1092[ 2 ] = fresh_wire_1098[ 0 ];
	assign fresh_wire_1092[ 3 ] = fresh_wire_1099[ 0 ];
	assign fresh_wire_1092[ 4 ] = fresh_wire_1100[ 0 ];
	assign fresh_wire_1092[ 5 ] = fresh_wire_1101[ 0 ];
	assign fresh_wire_1092[ 6 ] = fresh_wire_1102[ 0 ];
	assign fresh_wire_1092[ 7 ] = fresh_wire_1103[ 0 ];
	assign fresh_wire_1092[ 8 ] = fresh_wire_1104[ 0 ];
	assign fresh_wire_1093[ 0 ] = fresh_wire_435[ 0 ];
	assign fresh_wire_1093[ 1 ] = fresh_wire_435[ 1 ];
	assign fresh_wire_1093[ 2 ] = fresh_wire_435[ 2 ];
	assign fresh_wire_1093[ 3 ] = fresh_wire_435[ 3 ];
	assign fresh_wire_1093[ 4 ] = fresh_wire_435[ 4 ];
	assign fresh_wire_1093[ 5 ] = fresh_wire_435[ 5 ];
	assign fresh_wire_1093[ 6 ] = fresh_wire_435[ 6 ];
	assign fresh_wire_1093[ 7 ] = fresh_wire_435[ 7 ];
	assign fresh_wire_1093[ 8 ] = fresh_wire_435[ 8 ];
	assign fresh_wire_1095[ 0 ] = fresh_wire_1035[ 0 ];
	assign fresh_wire_1105[ 0 ] = fresh_wire_1109[ 0 ];
	assign fresh_wire_1105[ 1 ] = fresh_wire_1110[ 0 ];
	assign fresh_wire_1105[ 2 ] = fresh_wire_1111[ 0 ];
	assign fresh_wire_1105[ 3 ] = fresh_wire_1112[ 0 ];
	assign fresh_wire_1105[ 4 ] = fresh_wire_1113[ 0 ];
	assign fresh_wire_1105[ 5 ] = fresh_wire_1114[ 0 ];
	assign fresh_wire_1105[ 6 ] = fresh_wire_1115[ 0 ];
	assign fresh_wire_1105[ 7 ] = fresh_wire_1116[ 0 ];
	assign fresh_wire_1105[ 8 ] = fresh_wire_1117[ 0 ];
	assign fresh_wire_1106[ 0 ] = fresh_wire_1094[ 0 ];
	assign fresh_wire_1106[ 1 ] = fresh_wire_1094[ 1 ];
	assign fresh_wire_1106[ 2 ] = fresh_wire_1094[ 2 ];
	assign fresh_wire_1106[ 3 ] = fresh_wire_1094[ 3 ];
	assign fresh_wire_1106[ 4 ] = fresh_wire_1094[ 4 ];
	assign fresh_wire_1106[ 5 ] = fresh_wire_1094[ 5 ];
	assign fresh_wire_1106[ 6 ] = fresh_wire_1094[ 6 ];
	assign fresh_wire_1106[ 7 ] = fresh_wire_1094[ 7 ];
	assign fresh_wire_1106[ 8 ] = fresh_wire_1094[ 8 ];
	assign fresh_wire_1108[ 0 ] = fresh_wire_1032[ 0 ];
	assign fresh_wire_1118[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1119[ 0 ] = fresh_wire_435[ 0 ];
	assign fresh_wire_1119[ 1 ] = fresh_wire_435[ 1 ];
	assign fresh_wire_1119[ 2 ] = fresh_wire_435[ 2 ];
	assign fresh_wire_1119[ 3 ] = fresh_wire_435[ 3 ];
	assign fresh_wire_1119[ 4 ] = fresh_wire_435[ 4 ];
	assign fresh_wire_1119[ 5 ] = fresh_wire_435[ 5 ];
	assign fresh_wire_1119[ 6 ] = fresh_wire_435[ 6 ];
	assign fresh_wire_1119[ 7 ] = fresh_wire_435[ 7 ];
	assign fresh_wire_1119[ 8 ] = fresh_wire_435[ 8 ];
	assign fresh_wire_1121[ 0 ] = fresh_wire_1107[ 0 ];
	assign fresh_wire_1121[ 1 ] = fresh_wire_1107[ 1 ];
	assign fresh_wire_1121[ 2 ] = fresh_wire_1107[ 2 ];
	assign fresh_wire_1121[ 3 ] = fresh_wire_1107[ 3 ];
	assign fresh_wire_1121[ 4 ] = fresh_wire_1107[ 4 ];
	assign fresh_wire_1121[ 5 ] = fresh_wire_1107[ 5 ];
	assign fresh_wire_1121[ 6 ] = fresh_wire_1107[ 6 ];
	assign fresh_wire_1121[ 7 ] = fresh_wire_1107[ 7 ];
	assign fresh_wire_1121[ 8 ] = fresh_wire_1107[ 8 ];
	assign fresh_wire_1122[ 0 ] = fresh_wire_1074[ 0 ];
	assign fresh_wire_1122[ 1 ] = fresh_wire_1074[ 1 ];
	assign fresh_wire_1122[ 2 ] = fresh_wire_1074[ 2 ];
	assign fresh_wire_1122[ 3 ] = fresh_wire_1074[ 3 ];
	assign fresh_wire_1122[ 4 ] = fresh_wire_1074[ 4 ];
	assign fresh_wire_1122[ 5 ] = fresh_wire_1074[ 5 ];
	assign fresh_wire_1122[ 6 ] = fresh_wire_1074[ 6 ];
	assign fresh_wire_1122[ 7 ] = fresh_wire_1074[ 7 ];
	assign fresh_wire_1122[ 8 ] = fresh_wire_1074[ 8 ];
	assign fresh_wire_1122[ 9 ] = fresh_wire_1074[ 9 ];
	assign fresh_wire_1122[ 10 ] = fresh_wire_1074[ 10 ];
	assign fresh_wire_1122[ 11 ] = fresh_wire_1074[ 11 ];
	assign fresh_wire_1122[ 12 ] = fresh_wire_1074[ 12 ];
	assign fresh_wire_1122[ 13 ] = fresh_wire_1074[ 13 ];
	assign fresh_wire_1122[ 14 ] = fresh_wire_1074[ 14 ];
	assign fresh_wire_1122[ 15 ] = fresh_wire_1074[ 15 ];
	assign fresh_wire_1123[ 0 ] = fresh_wire_1050[ 0 ];
	assign fresh_wire_1124[ 0 ] = fresh_wire_96[ 0 ];
	assign fresh_wire_1124[ 1 ] = fresh_wire_94[ 0 ];
	assign fresh_wire_1124[ 2 ] = fresh_wire_92[ 0 ];
	assign fresh_wire_1124[ 3 ] = fresh_wire_90[ 0 ];
	assign fresh_wire_1124[ 4 ] = fresh_wire_88[ 0 ];
	assign fresh_wire_1124[ 5 ] = fresh_wire_86[ 0 ];
	assign fresh_wire_1124[ 6 ] = fresh_wire_114[ 0 ];
	assign fresh_wire_1124[ 7 ] = fresh_wire_112[ 0 ];
	assign fresh_wire_1124[ 8 ] = fresh_wire_110[ 0 ];
	assign fresh_wire_1124[ 9 ] = fresh_wire_108[ 0 ];
	assign fresh_wire_1124[ 10 ] = fresh_wire_106[ 0 ];
	assign fresh_wire_1124[ 11 ] = fresh_wire_104[ 0 ];
	assign fresh_wire_1124[ 12 ] = fresh_wire_102[ 0 ];
	assign fresh_wire_1124[ 13 ] = fresh_wire_100[ 0 ];
	assign fresh_wire_1124[ 14 ] = fresh_wire_98[ 0 ];
	assign fresh_wire_1124[ 15 ] = fresh_wire_84[ 0 ];
	assign fresh_wire_1124[ 16 ] = fresh_wire_1163[ 0 ];
	assign fresh_wire_1126[ 0 ] = fresh_wire_1125[ 0 ];
	assign fresh_wire_1126[ 1 ] = fresh_wire_1125[ 1 ];
	assign fresh_wire_1126[ 2 ] = fresh_wire_1125[ 2 ];
	assign fresh_wire_1126[ 3 ] = fresh_wire_1125[ 3 ];
	assign fresh_wire_1126[ 4 ] = fresh_wire_1125[ 4 ];
	assign fresh_wire_1126[ 5 ] = fresh_wire_1125[ 5 ];
	assign fresh_wire_1126[ 6 ] = fresh_wire_1125[ 6 ];
	assign fresh_wire_1126[ 7 ] = fresh_wire_1125[ 7 ];
	assign fresh_wire_1126[ 8 ] = fresh_wire_1125[ 8 ];
	assign fresh_wire_1126[ 9 ] = fresh_wire_1125[ 9 ];
	assign fresh_wire_1126[ 10 ] = fresh_wire_1125[ 10 ];
	assign fresh_wire_1126[ 11 ] = fresh_wire_1125[ 11 ];
	assign fresh_wire_1126[ 12 ] = fresh_wire_1125[ 12 ];
	assign fresh_wire_1126[ 13 ] = fresh_wire_1125[ 13 ];
	assign fresh_wire_1126[ 14 ] = fresh_wire_1125[ 14 ];
	assign fresh_wire_1126[ 15 ] = fresh_wire_1125[ 15 ];
	assign fresh_wire_1126[ 16 ] = fresh_wire_1125[ 16 ];
	assign fresh_wire_1126[ 17 ] = fresh_wire_1125[ 17 ];
	assign fresh_wire_1126[ 18 ] = fresh_wire_1125[ 18 ];
	assign fresh_wire_1126[ 19 ] = fresh_wire_1125[ 19 ];
	assign fresh_wire_1126[ 20 ] = fresh_wire_1125[ 20 ];
	assign fresh_wire_1126[ 21 ] = fresh_wire_1125[ 21 ];
	assign fresh_wire_1126[ 22 ] = fresh_wire_1125[ 22 ];
	assign fresh_wire_1126[ 23 ] = fresh_wire_1125[ 23 ];
	assign fresh_wire_1126[ 24 ] = fresh_wire_1125[ 24 ];
	assign fresh_wire_1126[ 25 ] = fresh_wire_1125[ 25 ];
	assign fresh_wire_1126[ 26 ] = fresh_wire_1125[ 26 ];
	assign fresh_wire_1126[ 27 ] = fresh_wire_1125[ 27 ];
	assign fresh_wire_1126[ 28 ] = fresh_wire_1125[ 28 ];
	assign fresh_wire_1126[ 29 ] = fresh_wire_1125[ 29 ];
	assign fresh_wire_1126[ 30 ] = fresh_wire_1125[ 30 ];
	assign fresh_wire_1126[ 31 ] = fresh_wire_1125[ 31 ];
	assign fresh_wire_1126[ 32 ] = fresh_wire_1125[ 32 ];
	assign fresh_wire_1126[ 33 ] = fresh_wire_1125[ 33 ];
	assign fresh_wire_1127[ 0 ] = fresh_wire_1164[ 0 ];
	assign fresh_wire_1127[ 1 ] = fresh_wire_1164[ 1 ];
	assign fresh_wire_1127[ 2 ] = fresh_wire_1164[ 2 ];
	assign fresh_wire_1127[ 3 ] = fresh_wire_1164[ 3 ];
	assign fresh_wire_1127[ 4 ] = fresh_wire_1164[ 4 ];
	assign fresh_wire_1127[ 5 ] = fresh_wire_1164[ 5 ];
	assign fresh_wire_1127[ 6 ] = fresh_wire_1164[ 6 ];
	assign fresh_wire_1127[ 7 ] = fresh_wire_1164[ 7 ];
	assign fresh_wire_1127[ 8 ] = fresh_wire_1164[ 8 ];
	assign fresh_wire_1127[ 9 ] = fresh_wire_1164[ 9 ];
	assign fresh_wire_1127[ 10 ] = fresh_wire_1164[ 10 ];
	assign fresh_wire_1127[ 11 ] = fresh_wire_1164[ 11 ];
	assign fresh_wire_1127[ 12 ] = fresh_wire_1164[ 12 ];
	assign fresh_wire_1127[ 13 ] = fresh_wire_1164[ 13 ];
	assign fresh_wire_1127[ 14 ] = fresh_wire_1164[ 14 ];
	assign fresh_wire_1127[ 15 ] = fresh_wire_1164[ 15 ];
	assign fresh_wire_1127[ 16 ] = fresh_wire_1164[ 16 ];
	assign fresh_wire_1127[ 17 ] = fresh_wire_1164[ 17 ];
	assign fresh_wire_1127[ 18 ] = fresh_wire_1164[ 18 ];
	assign fresh_wire_1127[ 19 ] = fresh_wire_1164[ 19 ];
	assign fresh_wire_1127[ 20 ] = fresh_wire_1164[ 20 ];
	assign fresh_wire_1127[ 21 ] = fresh_wire_1164[ 21 ];
	assign fresh_wire_1127[ 22 ] = fresh_wire_1164[ 22 ];
	assign fresh_wire_1127[ 23 ] = fresh_wire_1164[ 23 ];
	assign fresh_wire_1127[ 24 ] = fresh_wire_1164[ 24 ];
	assign fresh_wire_1127[ 25 ] = fresh_wire_1164[ 25 ];
	assign fresh_wire_1127[ 26 ] = fresh_wire_1164[ 26 ];
	assign fresh_wire_1127[ 27 ] = fresh_wire_1164[ 27 ];
	assign fresh_wire_1127[ 28 ] = fresh_wire_1164[ 28 ];
	assign fresh_wire_1127[ 29 ] = fresh_wire_1164[ 29 ];
	assign fresh_wire_1127[ 30 ] = fresh_wire_1164[ 30 ];
	assign fresh_wire_1127[ 31 ] = fresh_wire_1164[ 31 ];
	assign fresh_wire_1127[ 32 ] = fresh_wire_1164[ 32 ];
	assign fresh_wire_1127[ 33 ] = fresh_wire_1164[ 33 ];
	assign fresh_wire_1129[ 0 ] = fresh_wire_1141[ 0 ];
	assign fresh_wire_1129[ 1 ] = fresh_wire_1141[ 1 ];
	assign fresh_wire_1129[ 2 ] = fresh_wire_1141[ 2 ];
	assign fresh_wire_1129[ 3 ] = fresh_wire_1141[ 3 ];
	assign fresh_wire_1129[ 4 ] = fresh_wire_1141[ 4 ];
	assign fresh_wire_1129[ 5 ] = fresh_wire_1141[ 5 ];
	assign fresh_wire_1129[ 6 ] = fresh_wire_1141[ 6 ];
	assign fresh_wire_1129[ 7 ] = fresh_wire_1141[ 7 ];
	assign fresh_wire_1129[ 8 ] = fresh_wire_1141[ 8 ];
	assign fresh_wire_1129[ 9 ] = fresh_wire_1141[ 9 ];
	assign fresh_wire_1129[ 10 ] = fresh_wire_1141[ 10 ];
	assign fresh_wire_1129[ 11 ] = fresh_wire_1141[ 11 ];
	assign fresh_wire_1129[ 12 ] = fresh_wire_1141[ 12 ];
	assign fresh_wire_1129[ 13 ] = fresh_wire_1141[ 13 ];
	assign fresh_wire_1129[ 14 ] = fresh_wire_1141[ 14 ];
	assign fresh_wire_1129[ 15 ] = fresh_wire_1141[ 15 ];
	assign fresh_wire_1131[ 0 ] = fresh_wire_1130[ 0 ];
	assign fresh_wire_1131[ 1 ] = fresh_wire_1130[ 1 ];
	assign fresh_wire_1131[ 2 ] = fresh_wire_1130[ 2 ];
	assign fresh_wire_1131[ 3 ] = fresh_wire_1130[ 3 ];
	assign fresh_wire_1131[ 4 ] = fresh_wire_1130[ 4 ];
	assign fresh_wire_1131[ 5 ] = fresh_wire_1130[ 5 ];
	assign fresh_wire_1131[ 6 ] = fresh_wire_1130[ 6 ];
	assign fresh_wire_1131[ 7 ] = fresh_wire_1130[ 7 ];
	assign fresh_wire_1131[ 8 ] = fresh_wire_1130[ 8 ];
	assign fresh_wire_1131[ 9 ] = fresh_wire_1130[ 9 ];
	assign fresh_wire_1131[ 10 ] = fresh_wire_1130[ 10 ];
	assign fresh_wire_1131[ 11 ] = fresh_wire_1130[ 11 ];
	assign fresh_wire_1131[ 12 ] = fresh_wire_1130[ 12 ];
	assign fresh_wire_1131[ 13 ] = fresh_wire_1130[ 13 ];
	assign fresh_wire_1131[ 14 ] = fresh_wire_1130[ 14 ];
	assign fresh_wire_1131[ 15 ] = fresh_wire_1130[ 15 ];
	assign fresh_wire_1131[ 16 ] = fresh_wire_1130[ 16 ];
	assign fresh_wire_1132[ 0 ] = fresh_wire_1166[ 0 ];
	assign fresh_wire_1132[ 1 ] = fresh_wire_1166[ 1 ];
	assign fresh_wire_1132[ 2 ] = fresh_wire_1166[ 2 ];
	assign fresh_wire_1132[ 3 ] = fresh_wire_1166[ 3 ];
	assign fresh_wire_1132[ 4 ] = fresh_wire_1166[ 4 ];
	assign fresh_wire_1132[ 5 ] = fresh_wire_1166[ 5 ];
	assign fresh_wire_1132[ 6 ] = fresh_wire_1166[ 6 ];
	assign fresh_wire_1132[ 7 ] = fresh_wire_1166[ 7 ];
	assign fresh_wire_1132[ 8 ] = fresh_wire_1166[ 8 ];
	assign fresh_wire_1132[ 9 ] = fresh_wire_1166[ 9 ];
	assign fresh_wire_1132[ 10 ] = fresh_wire_1166[ 10 ];
	assign fresh_wire_1132[ 11 ] = fresh_wire_1166[ 11 ];
	assign fresh_wire_1132[ 12 ] = fresh_wire_1166[ 12 ];
	assign fresh_wire_1132[ 13 ] = fresh_wire_1166[ 13 ];
	assign fresh_wire_1132[ 14 ] = fresh_wire_1166[ 14 ];
	assign fresh_wire_1132[ 15 ] = fresh_wire_1166[ 15 ];
	assign fresh_wire_1132[ 16 ] = fresh_wire_1166[ 16 ];
	assign fresh_wire_1134[ 0 ] = fresh_wire_1133[ 0 ];
	assign fresh_wire_1134[ 1 ] = fresh_wire_1133[ 1 ];
	assign fresh_wire_1134[ 2 ] = fresh_wire_1133[ 2 ];
	assign fresh_wire_1134[ 3 ] = fresh_wire_1133[ 3 ];
	assign fresh_wire_1134[ 4 ] = fresh_wire_1133[ 4 ];
	assign fresh_wire_1134[ 5 ] = fresh_wire_1133[ 5 ];
	assign fresh_wire_1134[ 6 ] = fresh_wire_1133[ 6 ];
	assign fresh_wire_1134[ 7 ] = fresh_wire_1133[ 7 ];
	assign fresh_wire_1134[ 8 ] = fresh_wire_1133[ 8 ];
	assign fresh_wire_1134[ 9 ] = fresh_wire_1133[ 9 ];
	assign fresh_wire_1134[ 10 ] = fresh_wire_1133[ 10 ];
	assign fresh_wire_1134[ 11 ] = fresh_wire_1133[ 11 ];
	assign fresh_wire_1134[ 12 ] = fresh_wire_1133[ 12 ];
	assign fresh_wire_1134[ 13 ] = fresh_wire_1133[ 13 ];
	assign fresh_wire_1134[ 14 ] = fresh_wire_1133[ 14 ];
	assign fresh_wire_1134[ 15 ] = fresh_wire_1133[ 15 ];
	assign fresh_wire_1134[ 16 ] = fresh_wire_1133[ 16 ];
	assign fresh_wire_1135[ 0 ] = fresh_wire_1165[ 0 ];
	assign fresh_wire_1135[ 1 ] = fresh_wire_1165[ 1 ];
	assign fresh_wire_1135[ 2 ] = fresh_wire_1165[ 2 ];
	assign fresh_wire_1135[ 3 ] = fresh_wire_1165[ 3 ];
	assign fresh_wire_1135[ 4 ] = fresh_wire_1165[ 4 ];
	assign fresh_wire_1135[ 5 ] = fresh_wire_1165[ 5 ];
	assign fresh_wire_1135[ 6 ] = fresh_wire_1165[ 6 ];
	assign fresh_wire_1135[ 7 ] = fresh_wire_1165[ 7 ];
	assign fresh_wire_1135[ 8 ] = fresh_wire_1165[ 8 ];
	assign fresh_wire_1135[ 9 ] = fresh_wire_1165[ 9 ];
	assign fresh_wire_1135[ 10 ] = fresh_wire_1165[ 10 ];
	assign fresh_wire_1135[ 11 ] = fresh_wire_1165[ 11 ];
	assign fresh_wire_1135[ 12 ] = fresh_wire_1165[ 12 ];
	assign fresh_wire_1135[ 13 ] = fresh_wire_1165[ 13 ];
	assign fresh_wire_1135[ 14 ] = fresh_wire_1165[ 14 ];
	assign fresh_wire_1135[ 15 ] = fresh_wire_1165[ 15 ];
	assign fresh_wire_1135[ 16 ] = fresh_wire_1165[ 16 ];
	assign fresh_wire_1137[ 0 ] = fresh_wire_609[ 0 ];
	assign fresh_wire_1137[ 1 ] = fresh_wire_609[ 1 ];
	assign fresh_wire_1137[ 2 ] = fresh_wire_609[ 2 ];
	assign fresh_wire_1137[ 3 ] = fresh_wire_609[ 3 ];
	assign fresh_wire_1137[ 4 ] = fresh_wire_609[ 4 ];
	assign fresh_wire_1137[ 5 ] = fresh_wire_609[ 5 ];
	assign fresh_wire_1137[ 6 ] = fresh_wire_609[ 6 ];
	assign fresh_wire_1137[ 7 ] = fresh_wire_609[ 7 ];
	assign fresh_wire_1137[ 8 ] = fresh_wire_609[ 8 ];
	assign fresh_wire_1137[ 9 ] = fresh_wire_609[ 9 ];
	assign fresh_wire_1137[ 10 ] = fresh_wire_609[ 10 ];
	assign fresh_wire_1137[ 11 ] = fresh_wire_609[ 11 ];
	assign fresh_wire_1137[ 12 ] = fresh_wire_609[ 12 ];
	assign fresh_wire_1137[ 13 ] = fresh_wire_609[ 13 ];
	assign fresh_wire_1137[ 14 ] = fresh_wire_609[ 14 ];
	assign fresh_wire_1137[ 15 ] = fresh_wire_609[ 15 ];
	assign fresh_wire_1137[ 16 ] = fresh_wire_1167[ 0 ];
	assign fresh_wire_1139[ 0 ] = fresh_wire_1138[ 0 ];
	assign fresh_wire_1139[ 1 ] = fresh_wire_1138[ 1 ];
	assign fresh_wire_1139[ 2 ] = fresh_wire_1138[ 2 ];
	assign fresh_wire_1139[ 3 ] = fresh_wire_1138[ 3 ];
	assign fresh_wire_1139[ 4 ] = fresh_wire_1138[ 4 ];
	assign fresh_wire_1139[ 5 ] = fresh_wire_1138[ 5 ];
	assign fresh_wire_1139[ 6 ] = fresh_wire_1138[ 6 ];
	assign fresh_wire_1139[ 7 ] = fresh_wire_1138[ 7 ];
	assign fresh_wire_1139[ 8 ] = fresh_wire_1138[ 8 ];
	assign fresh_wire_1139[ 9 ] = fresh_wire_1138[ 9 ];
	assign fresh_wire_1139[ 10 ] = fresh_wire_1138[ 10 ];
	assign fresh_wire_1139[ 11 ] = fresh_wire_1138[ 11 ];
	assign fresh_wire_1139[ 12 ] = fresh_wire_1138[ 12 ];
	assign fresh_wire_1139[ 13 ] = fresh_wire_1138[ 13 ];
	assign fresh_wire_1139[ 14 ] = fresh_wire_1138[ 14 ];
	assign fresh_wire_1139[ 15 ] = fresh_wire_1138[ 15 ];
	assign fresh_wire_1139[ 16 ] = fresh_wire_1138[ 16 ];
	assign fresh_wire_1139[ 17 ] = fresh_wire_1138[ 17 ];
	assign fresh_wire_1139[ 18 ] = fresh_wire_1138[ 18 ];
	assign fresh_wire_1139[ 19 ] = fresh_wire_1138[ 19 ];
	assign fresh_wire_1139[ 20 ] = fresh_wire_1138[ 20 ];
	assign fresh_wire_1139[ 21 ] = fresh_wire_1138[ 21 ];
	assign fresh_wire_1139[ 22 ] = fresh_wire_1138[ 22 ];
	assign fresh_wire_1139[ 23 ] = fresh_wire_1138[ 23 ];
	assign fresh_wire_1139[ 24 ] = fresh_wire_1138[ 24 ];
	assign fresh_wire_1139[ 25 ] = fresh_wire_1138[ 25 ];
	assign fresh_wire_1139[ 26 ] = fresh_wire_1138[ 26 ];
	assign fresh_wire_1139[ 27 ] = fresh_wire_1138[ 27 ];
	assign fresh_wire_1139[ 28 ] = fresh_wire_1138[ 28 ];
	assign fresh_wire_1139[ 29 ] = fresh_wire_1138[ 29 ];
	assign fresh_wire_1139[ 30 ] = fresh_wire_1138[ 30 ];
	assign fresh_wire_1139[ 31 ] = fresh_wire_1138[ 31 ];
	assign fresh_wire_1139[ 32 ] = fresh_wire_1138[ 32 ];
	assign fresh_wire_1139[ 33 ] = fresh_wire_1138[ 33 ];
	assign fresh_wire_1140[ 0 ] = fresh_wire_1168[ 0 ];
	assign fresh_wire_1140[ 1 ] = fresh_wire_1168[ 1 ];
	assign fresh_wire_1140[ 2 ] = fresh_wire_1168[ 2 ];
	assign fresh_wire_1140[ 3 ] = fresh_wire_1168[ 3 ];
	assign fresh_wire_1140[ 4 ] = fresh_wire_1168[ 4 ];
	assign fresh_wire_1140[ 5 ] = fresh_wire_1168[ 5 ];
	assign fresh_wire_1140[ 6 ] = fresh_wire_1168[ 6 ];
	assign fresh_wire_1140[ 7 ] = fresh_wire_1168[ 7 ];
	assign fresh_wire_1140[ 8 ] = fresh_wire_1168[ 8 ];
	assign fresh_wire_1140[ 9 ] = fresh_wire_1168[ 9 ];
	assign fresh_wire_1140[ 10 ] = fresh_wire_1168[ 10 ];
	assign fresh_wire_1140[ 11 ] = fresh_wire_1168[ 11 ];
	assign fresh_wire_1140[ 12 ] = fresh_wire_1168[ 12 ];
	assign fresh_wire_1140[ 13 ] = fresh_wire_1168[ 13 ];
	assign fresh_wire_1140[ 14 ] = fresh_wire_1168[ 14 ];
	assign fresh_wire_1140[ 15 ] = fresh_wire_1168[ 15 ];
	assign fresh_wire_1140[ 16 ] = fresh_wire_1168[ 16 ];
	assign fresh_wire_1140[ 17 ] = fresh_wire_1168[ 17 ];
	assign fresh_wire_1140[ 18 ] = fresh_wire_1168[ 18 ];
	assign fresh_wire_1140[ 19 ] = fresh_wire_1168[ 19 ];
	assign fresh_wire_1140[ 20 ] = fresh_wire_1168[ 20 ];
	assign fresh_wire_1140[ 21 ] = fresh_wire_1168[ 21 ];
	assign fresh_wire_1140[ 22 ] = fresh_wire_1168[ 22 ];
	assign fresh_wire_1140[ 23 ] = fresh_wire_1168[ 23 ];
	assign fresh_wire_1140[ 24 ] = fresh_wire_1168[ 24 ];
	assign fresh_wire_1140[ 25 ] = fresh_wire_1168[ 25 ];
	assign fresh_wire_1140[ 26 ] = fresh_wire_1168[ 26 ];
	assign fresh_wire_1140[ 27 ] = fresh_wire_1168[ 27 ];
	assign fresh_wire_1140[ 28 ] = fresh_wire_1168[ 28 ];
	assign fresh_wire_1140[ 29 ] = fresh_wire_1168[ 29 ];
	assign fresh_wire_1140[ 30 ] = fresh_wire_1168[ 30 ];
	assign fresh_wire_1140[ 31 ] = fresh_wire_1168[ 31 ];
	assign fresh_wire_1140[ 32 ] = fresh_wire_1168[ 32 ];
	assign fresh_wire_1140[ 33 ] = fresh_wire_1168[ 33 ];
	assign fresh_wire_1142[ 0 ] = fresh_wire_1136[ 0 ];
	assign fresh_wire_1142[ 1 ] = fresh_wire_1136[ 1 ];
	assign fresh_wire_1142[ 2 ] = fresh_wire_1136[ 2 ];
	assign fresh_wire_1142[ 3 ] = fresh_wire_1136[ 3 ];
	assign fresh_wire_1142[ 4 ] = fresh_wire_1136[ 4 ];
	assign fresh_wire_1142[ 5 ] = fresh_wire_1136[ 5 ];
	assign fresh_wire_1142[ 6 ] = fresh_wire_1136[ 6 ];
	assign fresh_wire_1142[ 7 ] = fresh_wire_1136[ 7 ];
	assign fresh_wire_1142[ 8 ] = fresh_wire_1136[ 8 ];
	assign fresh_wire_1142[ 9 ] = fresh_wire_1136[ 9 ];
	assign fresh_wire_1142[ 10 ] = fresh_wire_1136[ 10 ];
	assign fresh_wire_1142[ 11 ] = fresh_wire_1136[ 11 ];
	assign fresh_wire_1142[ 12 ] = fresh_wire_1136[ 12 ];
	assign fresh_wire_1142[ 13 ] = fresh_wire_1136[ 13 ];
	assign fresh_wire_1142[ 14 ] = fresh_wire_1136[ 14 ];
	assign fresh_wire_1142[ 15 ] = fresh_wire_1136[ 15 ];
	assign fresh_wire_1144[ 0 ] = fresh_wire_1128[ 0 ];
	assign fresh_wire_1144[ 1 ] = fresh_wire_1128[ 1 ];
	assign fresh_wire_1144[ 2 ] = fresh_wire_1128[ 2 ];
	assign fresh_wire_1144[ 3 ] = fresh_wire_1128[ 3 ];
	assign fresh_wire_1144[ 4 ] = fresh_wire_1128[ 4 ];
	assign fresh_wire_1144[ 5 ] = fresh_wire_1128[ 5 ];
	assign fresh_wire_1144[ 6 ] = fresh_wire_1128[ 6 ];
	assign fresh_wire_1144[ 7 ] = fresh_wire_1128[ 7 ];
	assign fresh_wire_1144[ 8 ] = fresh_wire_1128[ 8 ];
	assign fresh_wire_1144[ 9 ] = fresh_wire_1128[ 9 ];
	assign fresh_wire_1144[ 10 ] = fresh_wire_1128[ 10 ];
	assign fresh_wire_1144[ 11 ] = fresh_wire_1128[ 11 ];
	assign fresh_wire_1144[ 12 ] = fresh_wire_1128[ 12 ];
	assign fresh_wire_1144[ 13 ] = fresh_wire_1128[ 13 ];
	assign fresh_wire_1144[ 14 ] = fresh_wire_1128[ 14 ];
	assign fresh_wire_1144[ 15 ] = fresh_wire_1128[ 15 ];
	assign fresh_wire_1146[ 0 ] = fresh_wire_1143[ 0 ];
	assign fresh_wire_1146[ 1 ] = fresh_wire_1143[ 1 ];
	assign fresh_wire_1146[ 2 ] = fresh_wire_1143[ 2 ];
	assign fresh_wire_1146[ 3 ] = fresh_wire_1143[ 3 ];
	assign fresh_wire_1146[ 4 ] = fresh_wire_1143[ 4 ];
	assign fresh_wire_1146[ 5 ] = fresh_wire_1143[ 5 ];
	assign fresh_wire_1146[ 6 ] = fresh_wire_1143[ 6 ];
	assign fresh_wire_1146[ 7 ] = fresh_wire_1143[ 7 ];
	assign fresh_wire_1146[ 8 ] = fresh_wire_1143[ 8 ];
	assign fresh_wire_1146[ 9 ] = fresh_wire_1143[ 9 ];
	assign fresh_wire_1146[ 10 ] = fresh_wire_1143[ 10 ];
	assign fresh_wire_1146[ 11 ] = fresh_wire_1143[ 11 ];
	assign fresh_wire_1146[ 12 ] = fresh_wire_1143[ 12 ];
	assign fresh_wire_1146[ 13 ] = fresh_wire_1143[ 13 ];
	assign fresh_wire_1146[ 14 ] = fresh_wire_1143[ 14 ];
	assign fresh_wire_1146[ 15 ] = fresh_wire_1143[ 15 ];
	assign fresh_wire_1146[ 16 ] = fresh_wire_1143[ 16 ];
	assign fresh_wire_1147[ 0 ] = fresh_wire_1145[ 0 ];
	assign fresh_wire_1147[ 1 ] = fresh_wire_1145[ 1 ];
	assign fresh_wire_1147[ 2 ] = fresh_wire_1145[ 2 ];
	assign fresh_wire_1147[ 3 ] = fresh_wire_1145[ 3 ];
	assign fresh_wire_1147[ 4 ] = fresh_wire_1145[ 4 ];
	assign fresh_wire_1147[ 5 ] = fresh_wire_1145[ 5 ];
	assign fresh_wire_1147[ 6 ] = fresh_wire_1145[ 6 ];
	assign fresh_wire_1147[ 7 ] = fresh_wire_1145[ 7 ];
	assign fresh_wire_1147[ 8 ] = fresh_wire_1145[ 8 ];
	assign fresh_wire_1147[ 9 ] = fresh_wire_1145[ 9 ];
	assign fresh_wire_1147[ 10 ] = fresh_wire_1145[ 10 ];
	assign fresh_wire_1147[ 11 ] = fresh_wire_1145[ 11 ];
	assign fresh_wire_1147[ 12 ] = fresh_wire_1145[ 12 ];
	assign fresh_wire_1147[ 13 ] = fresh_wire_1145[ 13 ];
	assign fresh_wire_1147[ 14 ] = fresh_wire_1145[ 14 ];
	assign fresh_wire_1147[ 15 ] = fresh_wire_1145[ 15 ];
	assign fresh_wire_1147[ 16 ] = fresh_wire_1145[ 16 ];
	assign fresh_wire_1149[ 0 ] = fresh_wire_1148[ 0 ];
	assign fresh_wire_1149[ 1 ] = fresh_wire_1148[ 1 ];
	assign fresh_wire_1149[ 2 ] = fresh_wire_1148[ 2 ];
	assign fresh_wire_1149[ 3 ] = fresh_wire_1148[ 3 ];
	assign fresh_wire_1149[ 4 ] = fresh_wire_1148[ 4 ];
	assign fresh_wire_1149[ 5 ] = fresh_wire_1148[ 5 ];
	assign fresh_wire_1149[ 6 ] = fresh_wire_1148[ 6 ];
	assign fresh_wire_1149[ 7 ] = fresh_wire_1148[ 7 ];
	assign fresh_wire_1149[ 8 ] = fresh_wire_1148[ 8 ];
	assign fresh_wire_1149[ 9 ] = fresh_wire_1148[ 9 ];
	assign fresh_wire_1149[ 10 ] = fresh_wire_1148[ 10 ];
	assign fresh_wire_1149[ 11 ] = fresh_wire_1148[ 11 ];
	assign fresh_wire_1149[ 12 ] = fresh_wire_1148[ 12 ];
	assign fresh_wire_1149[ 13 ] = fresh_wire_1148[ 13 ];
	assign fresh_wire_1149[ 14 ] = fresh_wire_1148[ 14 ];
	assign fresh_wire_1149[ 15 ] = fresh_wire_1148[ 15 ];
	assign fresh_wire_1149[ 16 ] = fresh_wire_1148[ 16 ];
	assign fresh_wire_1150[ 0 ] = fresh_wire_1174[ 0 ];
	assign fresh_wire_1150[ 1 ] = fresh_wire_1174[ 1 ];
	assign fresh_wire_1150[ 2 ] = fresh_wire_1174[ 2 ];
	assign fresh_wire_1150[ 3 ] = fresh_wire_1174[ 3 ];
	assign fresh_wire_1150[ 4 ] = fresh_wire_1174[ 4 ];
	assign fresh_wire_1150[ 5 ] = fresh_wire_1174[ 5 ];
	assign fresh_wire_1150[ 6 ] = fresh_wire_1174[ 6 ];
	assign fresh_wire_1150[ 7 ] = fresh_wire_1174[ 7 ];
	assign fresh_wire_1150[ 8 ] = fresh_wire_1174[ 8 ];
	assign fresh_wire_1150[ 9 ] = fresh_wire_1174[ 9 ];
	assign fresh_wire_1150[ 10 ] = fresh_wire_1174[ 10 ];
	assign fresh_wire_1150[ 11 ] = fresh_wire_1174[ 11 ];
	assign fresh_wire_1150[ 12 ] = fresh_wire_1174[ 12 ];
	assign fresh_wire_1150[ 13 ] = fresh_wire_1174[ 13 ];
	assign fresh_wire_1150[ 14 ] = fresh_wire_1174[ 14 ];
	assign fresh_wire_1150[ 15 ] = fresh_wire_1174[ 15 ];
	assign fresh_wire_1150[ 16 ] = fresh_wire_1174[ 16 ];
endmodule

