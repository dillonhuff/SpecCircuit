module CELL_TYPE_CONST #(parameter PARAM_WIDTH=1, parameter PARAM_INIT_VALUE=0) (output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT); assign PORT_ID_OUT = PARAM_INIT_VALUE;
endmodule

module CELL_TYPE_MUL #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT); assign PORT_ID_OUT = PORT_ID_IN0 * PORT_ID_IN1;
 endmodule

module CELL_TYPE_NOT #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT); assign PORT_ID_OUT = ~PORT_ID_IN;
 endmodule

module CELL_TYPE_ADD #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT);
   assign PORT_ID_OUT = PORT_ID_IN0 + PORT_ID_IN1;
 endmodule

module CELL_TYPE_SUB #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT);   assign PORT_ID_OUT = PORT_ID_IN0 - PORT_ID_IN1; endmodule

module CELL_TYPE_AND #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT);
   assign PORT_ID_OUT = PORT_ID_IN0 & PORT_ID_IN1;
endmodule

module CELL_TYPE_LSHR #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT);
   assign PORT_ID_OUT = PORT_ID_IN0 >> PORT_ID_IN1;
endmodule

module CELL_TYPE_ASHR #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT);
   assign PORT_ID_OUT = PORT_ID_IN0 >>> PORT_ID_IN1;
endmodule

module CELL_TYPE_XOR #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT);
   assign PORT_ID_OUT = PORT_ID_IN0 ^ PORT_ID_IN1;
endmodule

module CELL_TYPE_OR #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT);
   assign PORT_ID_OUT = PORT_ID_IN0 | PORT_ID_IN1;
endmodule

module CELL_TYPE_EQ #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [0 : 0] PORT_ID_OUT);
   assign PORT_ID_OUT = PORT_ID_IN0 == PORT_ID_IN1;
endmodule

module CELL_TYPE_NEQ #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [0 : 0] PORT_ID_OUT);
   assign PORT_ID_OUT = PORT_ID_IN0 != PORT_ID_IN1;
endmodule

module CELL_TYPE_ULT #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [0 : 0] PORT_ID_OUT); assign PORT_ID_OUT = PORT_ID_IN0 < PORT_ID_IN1;
 endmodule

module CELL_TYPE_UGE #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [0 : 0] PORT_ID_OUT); assign PORT_ID_OUT = PORT_ID_IN0 >= PORT_ID_IN1;
endmodule

 // CELL_TYPE_UGE
module CELL_TYPE_REG #(parameter PARAM_CLK_POSEDGE=1, parameter PARAM_INIT_VALUE=0, parameter PARAM_WIDTH=1)(input PORT_ID_CLK, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT);
   reg [PARAM_WIDTH - 1 : 0] data;
   initial begin
      data = PARAM_INIT_VALUE;
   end
   wire true_clk;
   assign true_clk = PARAM_CLK_POSEDGE ? PORT_ID_CLK : ~PORT_ID_CLK;
   always @(posedge true_clk) begin
      data <= PORT_ID_IN;
   end
   assign PORT_ID_OUT = data;
endmodule

module CELL_TYPE_REG_ARST #(parameter PARAM_CLK_POSEDGE=1, parameter PARAM_ARST_POSEDGE=1, parameter PARAM_INIT_VALUE=0, parameter PARAM_WIDTH=1)(input PORT_ID_ARST, input PORT_ID_CLK, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT);
   reg [PARAM_WIDTH - 1 : 0] data;
   initial begin
      data = PARAM_INIT_VALUE;
   end
   wire true_clk;
   assign true_clk = PARAM_CLK_POSEDGE ? PORT_ID_CLK : ~PORT_ID_CLK;
   wire true_rst;
   assign true_rst = PARAM_ARST_POSEDGE ? PORT_ID_ARST : ~PORT_ID_ARST;
   always @(posedge true_clk or posedge true_rst) begin
      if (true_rst) begin
         data <= PARAM_INIT_VALUE;
      end else begin
         data <= PORT_ID_IN;
      end
   end
   assign PORT_ID_OUT = data;
endmodule

 // CELL_TYPE_REG_ARST
module CELL_TYPE_MEM #(parameter PARAM_HAS_INIT=0, parameter PARAM_MEM_DEPTH=2, parameter PARAM_MEM_WIDTH=2)(input PORT_ID_CLK, input PORT_ID_WEN, input [$clog2(PARAM_MEM_DEPTH) - 1 : 0] PORT_ID_RADDR, input [$clog2(PARAM_MEM_DEPTH) - 1 : 0] PORT_ID_WADDR, input [PARAM_MEM_WIDTH - 1 : 0] PORT_ID_WDATA, output [PARAM_MEM_WIDTH - 1 : 0] PORT_ID_RDATA);
   reg [PARAM_MEM_WIDTH -  1 : 0] data_array [0 : PARAM_MEM_DEPTH - 1];
   always @(posedge PORT_ID_CLK) begin
      if (PORT_ID_WEN) begin
         data_array[PORT_ID_WADDR] = PORT_ID_WDATA;
      end
   end
   assign PORT_ID_RDATA = data_array[PORT_ID_RADDR];
endmodule

module CELL_TYPE_MUX #(parameter PARAM_WIDTH=1) (input PORT_ID_SEL, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT);
   assign PORT_ID_OUT = PORT_ID_SEL ? PORT_ID_IN1 : PORT_ID_IN0;
 endmodule

module CELL_TYPE_ORR #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN, output [0 : 0] PORT_ID_OUT); assign PORT_ID_OUT = |PORT_ID_IN;
 endmodule

module CELL_TYPE_ANDR #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN, output [0 : 0] PORT_ID_OUT); assign PORT_ID_OUT = &PORT_ID_IN;
 endmodule

module CELL_TYPE_PORT #(parameter PARAM_PORT_TYPE=0, parameter PARAM_OUT_WIDTH=1) (input [PARAM_OUT_WIDTH - 1 : 0] PORT_ID_IN, output [PARAM_OUT_WIDTH - 1 : 0] PORT_ID_OUT); assign PORT_ID_OUT = PORT_ID_IN;
 endmodule

module CELL_TYPE_ZEXT #(parameter PARAM_IN_WIDTH=1, parameter PARAM_OUT_WIDTH=1) (input [PARAM_IN_WIDTH - 1 : 0] PORT_ID_IN, output [PARAM_OUT_WIDTH - 1 : 0] PORT_ID_OUT); assign PORT_ID_OUT = {{(PARAM_OUT_WIDTH - PARAM_IN_WIDTH){1'b0}}, PORT_ID_IN};
 endmodule

module CELL_TYPE_SLICE #(parameter PARAM_WIDTH=1, parameter PARAM_LOW=1, parameter PARAM_HIGH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN, output [PARAM_HIGH - PARAM_LOW - 1 : 0] PORT_ID_OUT); assign PORT_ID_OUT = PORT_ID_IN[PARAM_HIGH:PARAM_LOW];
 endmodule

module CELL_TYPE_PASSTHROUGH #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT); assign PORT_ID_OUT = PORT_ID_IN;
 endmodule


module top(	output [0 : 0] aux_div_pad,
	input [0 : 0] clk_ext_in,
	input [0 : 0] clk_in,
	input [31 : 0] config_addr_in,
	input [31 : 0] config_data_in,
	input [0 : 0] ext_cki,
	input [0 : 0] ext_cki_jm,
	input [0 : 0] ext_ckib,
	input [0 : 0] ext_ckib_jm,
	input [0 : 0] ext_frefn,
	input [0 : 0] ext_frefn_jm,
	input [0 : 0] ext_frefp,
	input [0 : 0] ext_frefp_jm,
	output [0 : 0] ffeed_pad,
	output [0 : 0] fout_div_pad,
	output [0 : 0] fref_off_pad,
	output [0 : 0] frefn_out_jm,
	output [0 : 0] frefp_out_jm,
	output [12 : 0] lf_out,
	output [3 : 0] mdllout_pad,
	input [0 : 0] pad_S0_T0_in,
	output [0 : 0] pad_S0_T0_out,
	input [0 : 0] pad_S0_T10_in,
	output [0 : 0] pad_S0_T10_out,
	input [0 : 0] pad_S0_T11_in,
	output [0 : 0] pad_S0_T11_out,
	input [0 : 0] pad_S0_T12_in,
	output [0 : 0] pad_S0_T12_out,
	input [0 : 0] pad_S0_T13_in,
	output [0 : 0] pad_S0_T13_out,
	input [0 : 0] pad_S0_T14_in,
	output [0 : 0] pad_S0_T14_out,
	input [0 : 0] pad_S0_T15_in,
	output [0 : 0] pad_S0_T15_out,
	input [0 : 0] pad_S0_T1_in,
	output [0 : 0] pad_S0_T1_out,
	input [0 : 0] pad_S0_T2_in,
	output [0 : 0] pad_S0_T2_out,
	input [0 : 0] pad_S0_T3_in,
	output [0 : 0] pad_S0_T3_out,
	input [0 : 0] pad_S0_T4_in,
	output [0 : 0] pad_S0_T4_out,
	input [0 : 0] pad_S0_T5_in,
	output [0 : 0] pad_S0_T5_out,
	input [0 : 0] pad_S0_T6_in,
	output [0 : 0] pad_S0_T6_out,
	input [0 : 0] pad_S0_T7_in,
	output [0 : 0] pad_S0_T7_out,
	input [0 : 0] pad_S0_T8_in,
	output [0 : 0] pad_S0_T8_out,
	input [0 : 0] pad_S0_T9_in,
	output [0 : 0] pad_S0_T9_out,
	input [0 : 0] pad_S1_T0_in,
	output [0 : 0] pad_S1_T0_out,
	input [0 : 0] pad_S1_T10_in,
	output [0 : 0] pad_S1_T10_out,
	input [0 : 0] pad_S1_T11_in,
	output [0 : 0] pad_S1_T11_out,
	input [0 : 0] pad_S1_T12_in,
	output [0 : 0] pad_S1_T12_out,
	input [0 : 0] pad_S1_T13_in,
	output [0 : 0] pad_S1_T13_out,
	input [0 : 0] pad_S1_T14_in,
	output [0 : 0] pad_S1_T14_out,
	input [0 : 0] pad_S1_T15_in,
	output [0 : 0] pad_S1_T15_out,
	input [0 : 0] pad_S1_T1_in,
	output [0 : 0] pad_S1_T1_out,
	input [0 : 0] pad_S1_T2_in,
	output [0 : 0] pad_S1_T2_out,
	input [0 : 0] pad_S1_T3_in,
	output [0 : 0] pad_S1_T3_out,
	input [0 : 0] pad_S1_T4_in,
	output [0 : 0] pad_S1_T4_out,
	input [0 : 0] pad_S1_T5_in,
	output [0 : 0] pad_S1_T5_out,
	input [0 : 0] pad_S1_T6_in,
	output [0 : 0] pad_S1_T6_out,
	input [0 : 0] pad_S1_T7_in,
	output [0 : 0] pad_S1_T7_out,
	input [0 : 0] pad_S1_T8_in,
	output [0 : 0] pad_S1_T8_out,
	input [0 : 0] pad_S1_T9_in,
	output [0 : 0] pad_S1_T9_out,
	input [0 : 0] pad_S2_T0_in,
	output [0 : 0] pad_S2_T0_out,
	input [0 : 0] pad_S2_T10_in,
	output [0 : 0] pad_S2_T10_out,
	input [0 : 0] pad_S2_T11_in,
	output [0 : 0] pad_S2_T11_out,
	input [0 : 0] pad_S2_T12_in,
	output [0 : 0] pad_S2_T12_out,
	input [0 : 0] pad_S2_T13_in,
	output [0 : 0] pad_S2_T13_out,
	input [0 : 0] pad_S2_T14_in,
	output [0 : 0] pad_S2_T14_out,
	input [0 : 0] pad_S2_T15_in,
	output [0 : 0] pad_S2_T15_out,
	input [0 : 0] pad_S2_T1_in,
	output [0 : 0] pad_S2_T1_out,
	input [0 : 0] pad_S2_T2_in,
	output [0 : 0] pad_S2_T2_out,
	input [0 : 0] pad_S2_T3_in,
	output [0 : 0] pad_S2_T3_out,
	input [0 : 0] pad_S2_T4_in,
	output [0 : 0] pad_S2_T4_out,
	input [0 : 0] pad_S2_T5_in,
	output [0 : 0] pad_S2_T5_out,
	input [0 : 0] pad_S2_T6_in,
	output [0 : 0] pad_S2_T6_out,
	input [0 : 0] pad_S2_T7_in,
	output [0 : 0] pad_S2_T7_out,
	input [0 : 0] pad_S2_T8_in,
	output [0 : 0] pad_S2_T8_out,
	input [0 : 0] pad_S2_T9_in,
	output [0 : 0] pad_S2_T9_out,
	input [0 : 0] pad_S3_T0_in,
	output [0 : 0] pad_S3_T0_out,
	input [0 : 0] pad_S3_T10_in,
	output [0 : 0] pad_S3_T10_out,
	input [0 : 0] pad_S3_T11_in,
	output [0 : 0] pad_S3_T11_out,
	input [0 : 0] pad_S3_T12_in,
	output [0 : 0] pad_S3_T12_out,
	input [0 : 0] pad_S3_T13_in,
	output [0 : 0] pad_S3_T13_out,
	input [0 : 0] pad_S3_T14_in,
	output [0 : 0] pad_S3_T14_out,
	input [0 : 0] pad_S3_T15_in,
	output [0 : 0] pad_S3_T15_out,
	input [0 : 0] pad_S3_T1_in,
	output [0 : 0] pad_S3_T1_out,
	input [0 : 0] pad_S3_T2_in,
	output [0 : 0] pad_S3_T2_out,
	input [0 : 0] pad_S3_T3_in,
	output [0 : 0] pad_S3_T3_out,
	input [0 : 0] pad_S3_T4_in,
	output [0 : 0] pad_S3_T4_out,
	input [0 : 0] pad_S3_T5_in,
	output [0 : 0] pad_S3_T5_out,
	input [0 : 0] pad_S3_T6_in,
	output [0 : 0] pad_S3_T6_out,
	input [0 : 0] pad_S3_T7_in,
	output [0 : 0] pad_S3_T7_out,
	input [0 : 0] pad_S3_T8_in,
	output [0 : 0] pad_S3_T8_out,
	input [0 : 0] pad_S3_T9_in,
	output [0 : 0] pad_S3_T9_out,
	input [0 : 0] reset_in,
	input [0 : 0] tck,
	input [0 : 0] tdi,
	output [0 : 0] tdo,
	input [0 : 0] tms,
	input [0 : 0] trst_n);

	wire [0 : 0] fresh_wire_0;
	wire [0 : 0] fresh_wire_1;
	wire [0 : 0] fresh_wire_2;
	wire [31 : 0] fresh_wire_3;
	wire [31 : 0] fresh_wire_4;
	wire [0 : 0] fresh_wire_5;
	wire [0 : 0] fresh_wire_6;
	wire [0 : 0] fresh_wire_7;
	wire [0 : 0] fresh_wire_8;
	wire [0 : 0] fresh_wire_9;
	wire [0 : 0] fresh_wire_10;
	wire [0 : 0] fresh_wire_11;
	wire [0 : 0] fresh_wire_12;
	wire [0 : 0] fresh_wire_13;
	wire [0 : 0] fresh_wire_14;
	wire [0 : 0] fresh_wire_15;
	wire [0 : 0] fresh_wire_16;
	wire [0 : 0] fresh_wire_17;
	wire [12 : 0] fresh_wire_18;
	wire [3 : 0] fresh_wire_19;
	wire [0 : 0] fresh_wire_20;
	wire [0 : 0] fresh_wire_21;
	wire [0 : 0] fresh_wire_22;
	wire [0 : 0] fresh_wire_23;
	wire [0 : 0] fresh_wire_24;
	wire [0 : 0] fresh_wire_25;
	wire [0 : 0] fresh_wire_26;
	wire [0 : 0] fresh_wire_27;
	wire [0 : 0] fresh_wire_28;
	wire [0 : 0] fresh_wire_29;
	wire [0 : 0] fresh_wire_30;
	wire [0 : 0] fresh_wire_31;
	wire [0 : 0] fresh_wire_32;
	wire [0 : 0] fresh_wire_33;
	wire [0 : 0] fresh_wire_34;
	wire [0 : 0] fresh_wire_35;
	wire [0 : 0] fresh_wire_36;
	wire [0 : 0] fresh_wire_37;
	wire [0 : 0] fresh_wire_38;
	wire [0 : 0] fresh_wire_39;
	wire [0 : 0] fresh_wire_40;
	wire [0 : 0] fresh_wire_41;
	wire [0 : 0] fresh_wire_42;
	wire [0 : 0] fresh_wire_43;
	wire [0 : 0] fresh_wire_44;
	wire [0 : 0] fresh_wire_45;
	wire [0 : 0] fresh_wire_46;
	wire [0 : 0] fresh_wire_47;
	wire [0 : 0] fresh_wire_48;
	wire [0 : 0] fresh_wire_49;
	wire [0 : 0] fresh_wire_50;
	wire [0 : 0] fresh_wire_51;
	wire [0 : 0] fresh_wire_52;
	wire [0 : 0] fresh_wire_53;
	wire [0 : 0] fresh_wire_54;
	wire [0 : 0] fresh_wire_55;
	wire [0 : 0] fresh_wire_56;
	wire [0 : 0] fresh_wire_57;
	wire [0 : 0] fresh_wire_58;
	wire [0 : 0] fresh_wire_59;
	wire [0 : 0] fresh_wire_60;
	wire [0 : 0] fresh_wire_61;
	wire [0 : 0] fresh_wire_62;
	wire [0 : 0] fresh_wire_63;
	wire [0 : 0] fresh_wire_64;
	wire [0 : 0] fresh_wire_65;
	wire [0 : 0] fresh_wire_66;
	wire [0 : 0] fresh_wire_67;
	wire [0 : 0] fresh_wire_68;
	wire [0 : 0] fresh_wire_69;
	wire [0 : 0] fresh_wire_70;
	wire [0 : 0] fresh_wire_71;
	wire [0 : 0] fresh_wire_72;
	wire [0 : 0] fresh_wire_73;
	wire [0 : 0] fresh_wire_74;
	wire [0 : 0] fresh_wire_75;
	wire [0 : 0] fresh_wire_76;
	wire [0 : 0] fresh_wire_77;
	wire [0 : 0] fresh_wire_78;
	wire [0 : 0] fresh_wire_79;
	wire [0 : 0] fresh_wire_80;
	wire [0 : 0] fresh_wire_81;
	wire [0 : 0] fresh_wire_82;
	wire [0 : 0] fresh_wire_83;
	wire [0 : 0] fresh_wire_84;
	wire [0 : 0] fresh_wire_85;
	wire [0 : 0] fresh_wire_86;
	wire [0 : 0] fresh_wire_87;
	wire [0 : 0] fresh_wire_88;
	wire [0 : 0] fresh_wire_89;
	wire [0 : 0] fresh_wire_90;
	wire [0 : 0] fresh_wire_91;
	wire [0 : 0] fresh_wire_92;
	wire [0 : 0] fresh_wire_93;
	wire [0 : 0] fresh_wire_94;
	wire [0 : 0] fresh_wire_95;
	wire [0 : 0] fresh_wire_96;
	wire [0 : 0] fresh_wire_97;
	wire [0 : 0] fresh_wire_98;
	wire [0 : 0] fresh_wire_99;
	wire [0 : 0] fresh_wire_100;
	wire [0 : 0] fresh_wire_101;
	wire [0 : 0] fresh_wire_102;
	wire [0 : 0] fresh_wire_103;
	wire [0 : 0] fresh_wire_104;
	wire [0 : 0] fresh_wire_105;
	wire [0 : 0] fresh_wire_106;
	wire [0 : 0] fresh_wire_107;
	wire [0 : 0] fresh_wire_108;
	wire [0 : 0] fresh_wire_109;
	wire [0 : 0] fresh_wire_110;
	wire [0 : 0] fresh_wire_111;
	wire [0 : 0] fresh_wire_112;
	wire [0 : 0] fresh_wire_113;
	wire [0 : 0] fresh_wire_114;
	wire [0 : 0] fresh_wire_115;
	wire [0 : 0] fresh_wire_116;
	wire [0 : 0] fresh_wire_117;
	wire [0 : 0] fresh_wire_118;
	wire [0 : 0] fresh_wire_119;
	wire [0 : 0] fresh_wire_120;
	wire [0 : 0] fresh_wire_121;
	wire [0 : 0] fresh_wire_122;
	wire [0 : 0] fresh_wire_123;
	wire [0 : 0] fresh_wire_124;
	wire [0 : 0] fresh_wire_125;
	wire [0 : 0] fresh_wire_126;
	wire [0 : 0] fresh_wire_127;
	wire [0 : 0] fresh_wire_128;
	wire [0 : 0] fresh_wire_129;
	wire [0 : 0] fresh_wire_130;
	wire [0 : 0] fresh_wire_131;
	wire [0 : 0] fresh_wire_132;
	wire [0 : 0] fresh_wire_133;
	wire [0 : 0] fresh_wire_134;
	wire [0 : 0] fresh_wire_135;
	wire [0 : 0] fresh_wire_136;
	wire [0 : 0] fresh_wire_137;
	wire [0 : 0] fresh_wire_138;
	wire [0 : 0] fresh_wire_139;
	wire [0 : 0] fresh_wire_140;
	wire [0 : 0] fresh_wire_141;
	wire [0 : 0] fresh_wire_142;
	wire [0 : 0] fresh_wire_143;
	wire [0 : 0] fresh_wire_144;
	wire [0 : 0] fresh_wire_145;
	wire [0 : 0] fresh_wire_146;
	wire [0 : 0] fresh_wire_147;
	wire [0 : 0] fresh_wire_148;
	wire [0 : 0] fresh_wire_149;
	wire [0 : 0] fresh_wire_150;
	wire [0 : 0] fresh_wire_151;
	wire [0 : 0] fresh_wire_152;
	wire [0 : 0] fresh_wire_153;
	wire [12 : 0] fresh_wire_154;
	wire [0 : 0] fresh_wire_155;
	wire [0 : 0] fresh_wire_156;
	wire [0 : 0] fresh_wire_157;
	wire [0 : 0] fresh_wire_158;
	wire [0 : 0] fresh_wire_159;
	wire [0 : 0] fresh_wire_160;
	wire [0 : 0] fresh_wire_161;
	wire [0 : 0] fresh_wire_162;
	wire [0 : 0] fresh_wire_163;
	wire [15 : 0] fresh_wire_164;
	wire [15 : 0] fresh_wire_165;
	wire [15 : 0] fresh_wire_166;
	wire [1 : 0] fresh_wire_167;
	wire [15 : 0] fresh_wire_168;
	wire [15 : 0] fresh_wire_169;
	wire [15 : 0] fresh_wire_170;
	wire [15 : 0] fresh_wire_171;
	wire [15 : 0] fresh_wire_172;
	wire [31 : 0] fresh_wire_173;
	wire [31 : 0] fresh_wire_174;
	wire [31 : 0] fresh_wire_175;
	wire [31 : 0] fresh_wire_176;
	wire [15 : 0] fresh_wire_177;
	wire [31 : 0] fresh_wire_178;
	wire [31 : 0] fresh_wire_179;
	wire [31 : 0] fresh_wire_180;
	wire [31 : 0] fresh_wire_181;
	wire [15 : 0] fresh_wire_182;
	wire [31 : 0] fresh_wire_183;
	wire [31 : 0] fresh_wire_184;
	wire [31 : 0] fresh_wire_185;
	wire [31 : 0] fresh_wire_186;
	wire [15 : 0] fresh_wire_187;
	wire [15 : 0] fresh_wire_188;
	wire [15 : 0] fresh_wire_189;
	wire [15 : 0] fresh_wire_190;
	wire [15 : 0] fresh_wire_191;
	wire [15 : 0] fresh_wire_192;
	wire [15 : 0] fresh_wire_193;
	wire [15 : 0] fresh_wire_194;
	wire [15 : 0] fresh_wire_195;
	wire [15 : 0] fresh_wire_196;
	wire [15 : 0] fresh_wire_197;
	wire [15 : 0] fresh_wire_198;
	wire [0 : 0] fresh_wire_199;
	wire [0 : 0] fresh_wire_200;
	wire [0 : 0] fresh_wire_201;
	wire [1 : 0] fresh_wire_202;
	wire [1 : 0] fresh_wire_203;
	wire [0 : 0] fresh_wire_204;
	wire [1 : 0] fresh_wire_205;
	wire [1 : 0] fresh_wire_206;
	wire [0 : 0] fresh_wire_207;
	wire [1 : 0] fresh_wire_208;
	wire [1 : 0] fresh_wire_209;
	wire [0 : 0] fresh_wire_210;
	wire [15 : 0] fresh_wire_211;
	wire [15 : 0] fresh_wire_212;
	wire [0 : 0] fresh_wire_213;
	wire [0 : 0] fresh_wire_214;
	wire [0 : 0] fresh_wire_215;
	wire [0 : 0] fresh_wire_216;
	wire [0 : 0] fresh_wire_217;
	wire [0 : 0] fresh_wire_218;
	wire [0 : 0] fresh_wire_219;
	wire [0 : 0] fresh_wire_220;
	wire [0 : 0] fresh_wire_221;
	wire [0 : 0] fresh_wire_222;
	wire [0 : 0] fresh_wire_223;
	wire [0 : 0] fresh_wire_224;
	wire [0 : 0] fresh_wire_225;
	wire [1 : 0] fresh_wire_226;
	wire [1 : 0] fresh_wire_227;
	wire [0 : 0] fresh_wire_228;
	wire [0 : 0] fresh_wire_229;
	wire [0 : 0] fresh_wire_230;
	wire [0 : 0] fresh_wire_231;
	wire [0 : 0] fresh_wire_232;
	wire [0 : 0] fresh_wire_233;
	wire [0 : 0] fresh_wire_234;
	wire [1 : 0] fresh_wire_235;
	wire [1 : 0] fresh_wire_236;
	wire [0 : 0] fresh_wire_237;
	wire [0 : 0] fresh_wire_238;
	wire [0 : 0] fresh_wire_239;
	wire [0 : 0] fresh_wire_240;
	wire [0 : 0] fresh_wire_241;
	wire [0 : 0] fresh_wire_242;
	wire [0 : 0] fresh_wire_243;
	wire [1 : 0] fresh_wire_244;
	wire [1 : 0] fresh_wire_245;
	wire [0 : 0] fresh_wire_246;
	wire [1 : 0] fresh_wire_247;
	wire [1 : 0] fresh_wire_248;
	wire [0 : 0] fresh_wire_249;
	wire [15 : 0] fresh_wire_250;
	wire [15 : 0] fresh_wire_251;
	wire [0 : 0] fresh_wire_252;
	wire [0 : 0] fresh_wire_253;
	wire [0 : 0] fresh_wire_254;
	wire [0 : 0] fresh_wire_255;
	wire [0 : 0] fresh_wire_256;
	wire [0 : 0] fresh_wire_257;
	wire [0 : 0] fresh_wire_258;
	wire [15 : 0] fresh_wire_259;
	wire [15 : 0] fresh_wire_260;
	wire [0 : 0] fresh_wire_261;
	wire [15 : 0] fresh_wire_262;
	wire [15 : 0] fresh_wire_263;
	wire [0 : 0] fresh_wire_264;
	wire [15 : 0] fresh_wire_265;
	wire [15 : 0] fresh_wire_266;
	wire [0 : 0] fresh_wire_267;
	wire [0 : 0] fresh_wire_268;
	wire [0 : 0] fresh_wire_269;
	wire [0 : 0] fresh_wire_270;
	wire [0 : 0] fresh_wire_271;
	wire [0 : 0] fresh_wire_272;
	wire [0 : 0] fresh_wire_273;
	wire [0 : 0] fresh_wire_274;
	wire [0 : 0] fresh_wire_275;
	wire [0 : 0] fresh_wire_276;
	wire [0 : 0] fresh_wire_277;
	wire [0 : 0] fresh_wire_278;
	wire [0 : 0] fresh_wire_279;
	wire [0 : 0] fresh_wire_280;
	wire [0 : 0] fresh_wire_281;
	wire [0 : 0] fresh_wire_282;
	wire [0 : 0] fresh_wire_283;
	wire [0 : 0] fresh_wire_284;
	wire [0 : 0] fresh_wire_285;
	wire [0 : 0] fresh_wire_286;
	wire [0 : 0] fresh_wire_287;
	wire [0 : 0] fresh_wire_288;
	wire [0 : 0] fresh_wire_289;
	wire [0 : 0] fresh_wire_290;
	wire [0 : 0] fresh_wire_291;
	wire [0 : 0] fresh_wire_292;
	wire [0 : 0] fresh_wire_293;
	wire [0 : 0] fresh_wire_294;
	wire [0 : 0] fresh_wire_295;
	wire [0 : 0] fresh_wire_296;
	wire [0 : 0] fresh_wire_297;
	wire [0 : 0] fresh_wire_298;
	wire [0 : 0] fresh_wire_299;
	wire [0 : 0] fresh_wire_300;
	wire [0 : 0] fresh_wire_301;
	wire [0 : 0] fresh_wire_302;
	wire [0 : 0] fresh_wire_303;
	wire [0 : 0] fresh_wire_304;
	wire [0 : 0] fresh_wire_305;
	wire [0 : 0] fresh_wire_306;
	wire [0 : 0] fresh_wire_307;
	wire [0 : 0] fresh_wire_308;
	wire [0 : 0] fresh_wire_309;
	wire [0 : 0] fresh_wire_310;
	wire [0 : 0] fresh_wire_311;
	wire [0 : 0] fresh_wire_312;
	wire [0 : 0] fresh_wire_313;
	wire [0 : 0] fresh_wire_314;
	wire [0 : 0] fresh_wire_315;
	wire [0 : 0] fresh_wire_316;
	wire [0 : 0] fresh_wire_317;
	wire [0 : 0] fresh_wire_318;
	wire [0 : 0] fresh_wire_319;
	wire [0 : 0] fresh_wire_320;
	wire [0 : 0] fresh_wire_321;
	wire [0 : 0] fresh_wire_322;
	wire [0 : 0] fresh_wire_323;
	wire [0 : 0] fresh_wire_324;
	wire [0 : 0] fresh_wire_325;
	wire [0 : 0] fresh_wire_326;
	wire [0 : 0] fresh_wire_327;
	wire [0 : 0] fresh_wire_328;
	wire [0 : 0] fresh_wire_329;
	wire [0 : 0] fresh_wire_330;
	wire [0 : 0] fresh_wire_331;
	wire [0 : 0] fresh_wire_332;
	wire [0 : 0] fresh_wire_333;
	wire [0 : 0] fresh_wire_334;
	wire [0 : 0] fresh_wire_335;
	wire [0 : 0] fresh_wire_336;
	wire [0 : 0] fresh_wire_337;
	wire [0 : 0] fresh_wire_338;
	wire [0 : 0] fresh_wire_339;
	wire [0 : 0] fresh_wire_340;
	wire [0 : 0] fresh_wire_341;
	wire [0 : 0] fresh_wire_342;
	wire [0 : 0] fresh_wire_343;
	wire [0 : 0] fresh_wire_344;
	wire [0 : 0] fresh_wire_345;
	wire [0 : 0] fresh_wire_346;
	wire [0 : 0] fresh_wire_347;
	wire [0 : 0] fresh_wire_348;
	wire [0 : 0] fresh_wire_349;
	wire [0 : 0] fresh_wire_350;
	wire [0 : 0] fresh_wire_351;
	wire [0 : 0] fresh_wire_352;
	wire [0 : 0] fresh_wire_353;
	wire [0 : 0] fresh_wire_354;
	wire [0 : 0] fresh_wire_355;
	wire [0 : 0] fresh_wire_356;
	wire [0 : 0] fresh_wire_357;
	wire [0 : 0] fresh_wire_358;
	wire [0 : 0] fresh_wire_359;
	wire [0 : 0] fresh_wire_360;
	wire [15 : 0] fresh_wire_361;
	wire [15 : 0] fresh_wire_362;
	wire [0 : 0] fresh_wire_363;
	wire [15 : 0] fresh_wire_364;
	wire [15 : 0] fresh_wire_365;
	wire [0 : 0] fresh_wire_366;
	wire [0 : 0] fresh_wire_367;
	wire [0 : 0] fresh_wire_368;
	wire [0 : 0] fresh_wire_369;
	wire [0 : 0] fresh_wire_370;
	wire [0 : 0] fresh_wire_371;
	wire [1 : 0] fresh_wire_372;
	wire [1 : 0] fresh_wire_373;
	wire [0 : 0] fresh_wire_374;
	wire [1 : 0] fresh_wire_375;
	wire [1 : 0] fresh_wire_376;
	wire [0 : 0] fresh_wire_377;
	wire [15 : 0] fresh_wire_378;
	wire [15 : 0] fresh_wire_379;
	wire [0 : 0] fresh_wire_380;
	wire [0 : 0] fresh_wire_381;
	wire [0 : 0] fresh_wire_382;
	wire [0 : 0] fresh_wire_383;
	wire [0 : 0] fresh_wire_384;
	wire [0 : 0] fresh_wire_385;
	wire [0 : 0] fresh_wire_386;
	wire [0 : 0] fresh_wire_387;
	wire [0 : 0] fresh_wire_388;
	wire [0 : 0] fresh_wire_389;
	wire [0 : 0] fresh_wire_390;
	wire [0 : 0] fresh_wire_391;
	wire [0 : 0] fresh_wire_392;
	wire [0 : 0] fresh_wire_393;
	wire [0 : 0] fresh_wire_394;
	wire [0 : 0] fresh_wire_395;
	wire [0 : 0] fresh_wire_396;
	wire [0 : 0] fresh_wire_397;
	wire [0 : 0] fresh_wire_398;
	wire [0 : 0] fresh_wire_399;
	wire [0 : 0] fresh_wire_400;
	wire [1 : 0] fresh_wire_401;
	wire [1 : 0] fresh_wire_402;
	wire [0 : 0] fresh_wire_403;
	wire [0 : 0] fresh_wire_404;
	wire [15 : 0] fresh_wire_405;
	wire [15 : 0] fresh_wire_406;
	wire [0 : 0] fresh_wire_407;
	wire [0 : 0] fresh_wire_408;
	wire [15 : 0] fresh_wire_409;
	wire [15 : 0] fresh_wire_410;
	wire [0 : 0] fresh_wire_411;
	wire [0 : 0] fresh_wire_412;
	wire [15 : 0] fresh_wire_413;
	wire [15 : 0] fresh_wire_414;
	wire [0 : 0] fresh_wire_415;
	wire [0 : 0] fresh_wire_416;
	wire [15 : 0] fresh_wire_417;
	wire [15 : 0] fresh_wire_418;
	wire [0 : 0] fresh_wire_419;
	wire [0 : 0] fresh_wire_420;
	wire [0 : 0] fresh_wire_421;
	wire [0 : 0] fresh_wire_422;
	wire [0 : 0] fresh_wire_423;
	wire [0 : 0] fresh_wire_424;
	wire [0 : 0] fresh_wire_425;
	wire [0 : 0] fresh_wire_426;
	wire [0 : 0] fresh_wire_427;
	wire [0 : 0] fresh_wire_428;
	wire [0 : 0] fresh_wire_429;
	wire [0 : 0] fresh_wire_430;
	wire [0 : 0] fresh_wire_431;
	wire [0 : 0] fresh_wire_432;
	wire [15 : 0] fresh_wire_433;
	wire [15 : 0] fresh_wire_434;
	wire [15 : 0] fresh_wire_435;
	wire [0 : 0] fresh_wire_436;
	wire [0 : 0] fresh_wire_437;
	wire [0 : 0] fresh_wire_438;
	wire [0 : 0] fresh_wire_439;
	wire [0 : 0] fresh_wire_440;
	wire [0 : 0] fresh_wire_441;
	wire [0 : 0] fresh_wire_442;
	wire [0 : 0] fresh_wire_443;
	wire [0 : 0] fresh_wire_444;
	wire [0 : 0] fresh_wire_445;
	wire [0 : 0] fresh_wire_446;
	wire [0 : 0] fresh_wire_447;
	wire [0 : 0] fresh_wire_448;
	wire [0 : 0] fresh_wire_449;
	wire [0 : 0] fresh_wire_450;
	wire [0 : 0] fresh_wire_451;
	wire [0 : 0] fresh_wire_452;
	wire [0 : 0] fresh_wire_453;
	wire [0 : 0] fresh_wire_454;
	wire [0 : 0] fresh_wire_455;
	wire [0 : 0] fresh_wire_456;
	wire [15 : 0] fresh_wire_457;
	wire [15 : 0] fresh_wire_458;
	wire [15 : 0] fresh_wire_459;
	wire [0 : 0] fresh_wire_460;
	wire [15 : 0] fresh_wire_461;
	wire [15 : 0] fresh_wire_462;
	wire [15 : 0] fresh_wire_463;
	wire [0 : 0] fresh_wire_464;
	wire [15 : 0] fresh_wire_465;
	wire [15 : 0] fresh_wire_466;
	wire [15 : 0] fresh_wire_467;
	wire [0 : 0] fresh_wire_468;
	wire [15 : 0] fresh_wire_469;
	wire [15 : 0] fresh_wire_470;
	wire [15 : 0] fresh_wire_471;
	wire [0 : 0] fresh_wire_472;
	wire [1 : 0] fresh_wire_473;
	wire [1 : 0] fresh_wire_474;
	wire [1 : 0] fresh_wire_475;
	wire [0 : 0] fresh_wire_476;
	wire [1 : 0] fresh_wire_477;
	wire [1 : 0] fresh_wire_478;
	wire [1 : 0] fresh_wire_479;
	wire [0 : 0] fresh_wire_480;
	wire [1 : 0] fresh_wire_481;
	wire [1 : 0] fresh_wire_482;
	wire [1 : 0] fresh_wire_483;
	wire [0 : 0] fresh_wire_484;
	wire [1 : 0] fresh_wire_485;
	wire [1 : 0] fresh_wire_486;
	wire [1 : 0] fresh_wire_487;
	wire [0 : 0] fresh_wire_488;
	wire [1 : 0] fresh_wire_489;
	wire [1 : 0] fresh_wire_490;
	wire [1 : 0] fresh_wire_491;
	wire [0 : 0] fresh_wire_492;
	wire [1 : 0] fresh_wire_493;
	wire [1 : 0] fresh_wire_494;
	wire [1 : 0] fresh_wire_495;
	wire [0 : 0] fresh_wire_496;
	wire [0 : 0] fresh_wire_497;
	wire [0 : 0] fresh_wire_498;
	wire [0 : 0] fresh_wire_499;
	wire [0 : 0] fresh_wire_500;
	wire [0 : 0] fresh_wire_501;
	wire [0 : 0] fresh_wire_502;
	wire [0 : 0] fresh_wire_503;
	wire [0 : 0] fresh_wire_504;
	wire [0 : 0] fresh_wire_505;
	wire [0 : 0] fresh_wire_506;
	wire [0 : 0] fresh_wire_507;
	wire [0 : 0] fresh_wire_508;
	wire [0 : 0] fresh_wire_509;
	wire [0 : 0] fresh_wire_510;
	wire [0 : 0] fresh_wire_511;
	wire [0 : 0] fresh_wire_512;
	wire [0 : 0] fresh_wire_513;
	wire [0 : 0] fresh_wire_514;
	wire [0 : 0] fresh_wire_515;
	wire [0 : 0] fresh_wire_516;
	wire [0 : 0] fresh_wire_517;
	wire [0 : 0] fresh_wire_518;
	wire [0 : 0] fresh_wire_519;
	wire [0 : 0] fresh_wire_520;
	wire [0 : 0] fresh_wire_521;
	wire [0 : 0] fresh_wire_522;
	wire [0 : 0] fresh_wire_523;
	wire [0 : 0] fresh_wire_524;
	wire [0 : 0] fresh_wire_525;
	wire [0 : 0] fresh_wire_526;
	wire [0 : 0] fresh_wire_527;
	wire [0 : 0] fresh_wire_528;
	wire [0 : 0] fresh_wire_529;
	wire [0 : 0] fresh_wire_530;
	wire [0 : 0] fresh_wire_531;
	wire [0 : 0] fresh_wire_532;
	wire [0 : 0] fresh_wire_533;
	wire [0 : 0] fresh_wire_534;
	wire [0 : 0] fresh_wire_535;
	wire [0 : 0] fresh_wire_536;
	wire [15 : 0] fresh_wire_537;
	wire [15 : 0] fresh_wire_538;
	wire [15 : 0] fresh_wire_539;
	wire [0 : 0] fresh_wire_540;
	wire [15 : 0] fresh_wire_541;
	wire [15 : 0] fresh_wire_542;
	wire [15 : 0] fresh_wire_543;
	wire [0 : 0] fresh_wire_544;
	wire [15 : 0] fresh_wire_545;
	wire [15 : 0] fresh_wire_546;
	wire [15 : 0] fresh_wire_547;
	wire [0 : 0] fresh_wire_548;
	wire [15 : 0] fresh_wire_549;
	wire [15 : 0] fresh_wire_550;
	wire [15 : 0] fresh_wire_551;
	wire [0 : 0] fresh_wire_552;
	wire [15 : 0] fresh_wire_553;
	wire [15 : 0] fresh_wire_554;
	wire [15 : 0] fresh_wire_555;
	wire [0 : 0] fresh_wire_556;
	wire [15 : 0] fresh_wire_557;
	wire [15 : 0] fresh_wire_558;
	wire [15 : 0] fresh_wire_559;
	wire [0 : 0] fresh_wire_560;
	wire [15 : 0] fresh_wire_561;
	wire [15 : 0] fresh_wire_562;
	wire [15 : 0] fresh_wire_563;
	wire [0 : 0] fresh_wire_564;
	wire [15 : 0] fresh_wire_565;
	wire [15 : 0] fresh_wire_566;
	wire [15 : 0] fresh_wire_567;
	wire [0 : 0] fresh_wire_568;
	wire [15 : 0] fresh_wire_569;
	wire [15 : 0] fresh_wire_570;
	wire [15 : 0] fresh_wire_571;
	wire [0 : 0] fresh_wire_572;
	wire [0 : 0] fresh_wire_573;
	wire [0 : 0] fresh_wire_574;
	wire [0 : 0] fresh_wire_575;
	wire [0 : 0] fresh_wire_576;
	wire [0 : 0] fresh_wire_577;
	wire [0 : 0] fresh_wire_578;
	wire [0 : 0] fresh_wire_579;
	wire [0 : 0] fresh_wire_580;
	wire [0 : 0] fresh_wire_581;
	wire [0 : 0] fresh_wire_582;
	wire [0 : 0] fresh_wire_583;
	wire [0 : 0] fresh_wire_584;
	wire [0 : 0] fresh_wire_585;
	wire [0 : 0] fresh_wire_586;
	wire [0 : 0] fresh_wire_587;
	wire [0 : 0] fresh_wire_588;
	wire [0 : 0] fresh_wire_589;
	wire [0 : 0] fresh_wire_590;
	wire [0 : 0] fresh_wire_591;
	wire [0 : 0] fresh_wire_592;
	wire [15 : 0] fresh_wire_593;
	wire [31 : 0] fresh_wire_594;
	wire [31 : 0] fresh_wire_595;
	wire [31 : 0] fresh_wire_596;
	wire [31 : 0] fresh_wire_597;
	wire [31 : 0] fresh_wire_598;
	wire [31 : 0] fresh_wire_599;
	wire [31 : 0] fresh_wire_600;
	wire [0 : 0] fresh_wire_601;
	wire [15 : 0] fresh_wire_602;
	wire [15 : 0] fresh_wire_603;
	wire [15 : 0] fresh_wire_604;
	wire [0 : 0] fresh_wire_605;
	wire [0 : 0] fresh_wire_606;
	wire [15 : 0] fresh_wire_607;
	wire [15 : 0] fresh_wire_608;
	wire [15 : 0] fresh_wire_609;
	wire [0 : 0] fresh_wire_610;
	wire [1 : 0] fresh_wire_611;
	wire [1 : 0] fresh_wire_612;
	wire [1 : 0] fresh_wire_613;
	wire [0 : 0] fresh_wire_614;
	wire [0 : 0] fresh_wire_615;
	wire [0 : 0] fresh_wire_616;
	wire [0 : 0] fresh_wire_617;
	wire [0 : 0] fresh_wire_618;
	wire [0 : 0] fresh_wire_619;
	wire [0 : 0] fresh_wire_620;
	wire [0 : 0] fresh_wire_621;
	wire [0 : 0] fresh_wire_622;
	wire [1 : 0] fresh_wire_623;
	wire [1 : 0] fresh_wire_624;
	wire [0 : 0] fresh_wire_625;
	wire [1 : 0] fresh_wire_626;
	wire [1 : 0] fresh_wire_627;
	wire [0 : 0] fresh_wire_628;
	wire [0 : 0] fresh_wire_629;
	wire [0 : 0] fresh_wire_630;
	wire [0 : 0] fresh_wire_631;
	wire [1 : 0] fresh_wire_632;
	wire [1 : 0] fresh_wire_633;
	wire [0 : 0] fresh_wire_634;
	wire [1 : 0] fresh_wire_635;
	wire [1 : 0] fresh_wire_636;
	wire [0 : 0] fresh_wire_637;
	wire [0 : 0] fresh_wire_638;
	wire [0 : 0] fresh_wire_639;
	wire [0 : 0] fresh_wire_640;
	wire [0 : 0] fresh_wire_641;
	wire [0 : 0] fresh_wire_642;
	wire [0 : 0] fresh_wire_643;
	wire [0 : 0] fresh_wire_644;
	wire [0 : 0] fresh_wire_645;
	wire [0 : 0] fresh_wire_646;
	wire [0 : 0] fresh_wire_647;
	wire [0 : 0] fresh_wire_648;
	wire [0 : 0] fresh_wire_649;
	wire [0 : 0] fresh_wire_650;
	wire [0 : 0] fresh_wire_651;
	wire [0 : 0] fresh_wire_652;
	wire [0 : 0] fresh_wire_653;
	wire [0 : 0] fresh_wire_654;
	wire [0 : 0] fresh_wire_655;
	wire [0 : 0] fresh_wire_656;
	wire [0 : 0] fresh_wire_657;
	wire [0 : 0] fresh_wire_658;
	wire [0 : 0] fresh_wire_659;
	wire [0 : 0] fresh_wire_660;
	wire [0 : 0] fresh_wire_661;
	wire [0 : 0] fresh_wire_662;
	wire [0 : 0] fresh_wire_663;
	wire [0 : 0] fresh_wire_664;
	wire [1 : 0] fresh_wire_665;
	wire [1 : 0] fresh_wire_666;
	wire [0 : 0] fresh_wire_667;
	wire [0 : 0] fresh_wire_668;
	wire [47 : 0] fresh_wire_669;
	wire [47 : 0] fresh_wire_670;
	wire [0 : 0] fresh_wire_671;
	wire [0 : 0] fresh_wire_672;
	wire [0 : 0] fresh_wire_673;
	wire [0 : 0] fresh_wire_674;
	wire [0 : 0] fresh_wire_675;
	wire [0 : 0] fresh_wire_676;
	wire [0 : 0] fresh_wire_677;
	wire [0 : 0] fresh_wire_678;
	wire [0 : 0] fresh_wire_679;
	wire [1 : 0] fresh_wire_680;
	wire [1 : 0] fresh_wire_681;
	wire [1 : 0] fresh_wire_682;
	wire [0 : 0] fresh_wire_683;
	wire [1 : 0] fresh_wire_684;
	wire [1 : 0] fresh_wire_685;
	wire [1 : 0] fresh_wire_686;
	wire [0 : 0] fresh_wire_687;
	wire [31 : 0] fresh_wire_688;
	wire [31 : 0] fresh_wire_689;
	wire [31 : 0] fresh_wire_690;
	wire [0 : 0] fresh_wire_691;
	wire [31 : 0] fresh_wire_692;
	wire [31 : 0] fresh_wire_693;
	wire [31 : 0] fresh_wire_694;
	wire [0 : 0] fresh_wire_695;
	wire [31 : 0] fresh_wire_696;
	wire [31 : 0] fresh_wire_697;
	wire [31 : 0] fresh_wire_698;
	wire [0 : 0] fresh_wire_699;
	wire [31 : 0] fresh_wire_700;
	wire [31 : 0] fresh_wire_701;
	wire [31 : 0] fresh_wire_702;
	wire [0 : 0] fresh_wire_703;
	wire [31 : 0] fresh_wire_704;
	wire [31 : 0] fresh_wire_705;
	wire [31 : 0] fresh_wire_706;
	wire [0 : 0] fresh_wire_707;
	wire [31 : 0] fresh_wire_708;
	wire [31 : 0] fresh_wire_709;
	wire [31 : 0] fresh_wire_710;
	wire [0 : 0] fresh_wire_711;
	wire [31 : 0] fresh_wire_712;
	wire [31 : 0] fresh_wire_713;
	wire [31 : 0] fresh_wire_714;
	wire [0 : 0] fresh_wire_715;
	wire [1 : 0] fresh_wire_716;
	wire [1 : 0] fresh_wire_717;
	wire [1 : 0] fresh_wire_718;
	wire [0 : 0] fresh_wire_719;
	wire [1 : 0] fresh_wire_720;
	wire [1 : 0] fresh_wire_721;
	wire [1 : 0] fresh_wire_722;
	wire [1 : 0] fresh_wire_723;
	wire [1 : 0] fresh_wire_724;
	wire [1 : 0] fresh_wire_725;
	wire [0 : 0] fresh_wire_726;
	wire [0 : 0] fresh_wire_727;
	wire [0 : 0] fresh_wire_728;
	wire [0 : 0] fresh_wire_729;
	wire [0 : 0] fresh_wire_730;
	wire [0 : 0] fresh_wire_731;
	wire [0 : 0] fresh_wire_732;
	wire [0 : 0] fresh_wire_733;
	wire [0 : 0] fresh_wire_734;
	wire [0 : 0] fresh_wire_735;
	wire [0 : 0] fresh_wire_736;
	wire [0 : 0] fresh_wire_737;
	wire [0 : 0] fresh_wire_738;
	wire [0 : 0] fresh_wire_739;
	wire [0 : 0] fresh_wire_740;
	wire [0 : 0] fresh_wire_741;
	wire [0 : 0] fresh_wire_742;
	wire [0 : 0] fresh_wire_743;
	wire [1 : 0] fresh_wire_744;
	wire [1 : 0] fresh_wire_745;
	wire [0 : 0] fresh_wire_746;
	wire [1 : 0] fresh_wire_747;
	wire [1 : 0] fresh_wire_748;
	wire [0 : 0] fresh_wire_749;
	wire [1 : 0] fresh_wire_750;
	wire [1 : 0] fresh_wire_751;
	wire [0 : 0] fresh_wire_752;
	wire [1 : 0] fresh_wire_753;
	wire [1 : 0] fresh_wire_754;
	wire [0 : 0] fresh_wire_755;
	wire [1 : 0] fresh_wire_756;
	wire [1 : 0] fresh_wire_757;
	wire [0 : 0] fresh_wire_758;
	wire [0 : 0] fresh_wire_759;
	wire [0 : 0] fresh_wire_760;
	wire [0 : 0] fresh_wire_761;
	wire [0 : 0] fresh_wire_762;
	wire [0 : 0] fresh_wire_763;
	wire [0 : 0] fresh_wire_764;
	wire [0 : 0] fresh_wire_765;
	wire [0 : 0] fresh_wire_766;
	wire [0 : 0] fresh_wire_767;
	wire [0 : 0] fresh_wire_768;
	wire [0 : 0] fresh_wire_769;
	wire [0 : 0] fresh_wire_770;
	wire [0 : 0] fresh_wire_771;
	wire [0 : 0] fresh_wire_772;
	wire [0 : 0] fresh_wire_773;
	wire [0 : 0] fresh_wire_774;
	wire [0 : 0] fresh_wire_775;
	wire [0 : 0] fresh_wire_776;
	wire [0 : 0] fresh_wire_777;
	wire [0 : 0] fresh_wire_778;
	wire [0 : 0] fresh_wire_779;
	wire [0 : 0] fresh_wire_780;
	wire [0 : 0] fresh_wire_781;
	wire [0 : 0] fresh_wire_782;
	wire [0 : 0] fresh_wire_783;
	wire [0 : 0] fresh_wire_784;
	wire [0 : 0] fresh_wire_785;
	wire [0 : 0] fresh_wire_786;
	wire [0 : 0] fresh_wire_787;
	wire [0 : 0] fresh_wire_788;
	wire [0 : 0] fresh_wire_789;
	wire [0 : 0] fresh_wire_790;
	wire [0 : 0] fresh_wire_791;
	wire [0 : 0] fresh_wire_792;
	wire [0 : 0] fresh_wire_793;
	wire [0 : 0] fresh_wire_794;
	wire [0 : 0] fresh_wire_795;
	wire [0 : 0] fresh_wire_796;
	wire [0 : 0] fresh_wire_797;
	wire [0 : 0] fresh_wire_798;
	wire [0 : 0] fresh_wire_799;
	wire [0 : 0] fresh_wire_800;
	wire [0 : 0] fresh_wire_801;
	wire [0 : 0] fresh_wire_802;
	wire [0 : 0] fresh_wire_803;
	wire [0 : 0] fresh_wire_804;
	wire [0 : 0] fresh_wire_805;
	wire [0 : 0] fresh_wire_806;
	wire [0 : 0] fresh_wire_807;
	wire [0 : 0] fresh_wire_808;
	wire [0 : 0] fresh_wire_809;
	wire [0 : 0] fresh_wire_810;
	wire [0 : 0] fresh_wire_811;
	wire [0 : 0] fresh_wire_812;
	wire [0 : 0] fresh_wire_813;
	wire [0 : 0] fresh_wire_814;
	wire [0 : 0] fresh_wire_815;
	wire [0 : 0] fresh_wire_816;
	wire [0 : 0] fresh_wire_817;
	wire [0 : 0] fresh_wire_818;
	wire [0 : 0] fresh_wire_819;
	wire [0 : 0] fresh_wire_820;
	wire [0 : 0] fresh_wire_821;
	wire [0 : 0] fresh_wire_822;
	wire [0 : 0] fresh_wire_823;
	wire [0 : 0] fresh_wire_824;
	wire [0 : 0] fresh_wire_825;
	wire [0 : 0] fresh_wire_826;
	wire [0 : 0] fresh_wire_827;
	wire [0 : 0] fresh_wire_828;
	wire [0 : 0] fresh_wire_829;
	wire [0 : 0] fresh_wire_830;
	wire [0 : 0] fresh_wire_831;
	wire [0 : 0] fresh_wire_832;
	wire [0 : 0] fresh_wire_833;
	wire [0 : 0] fresh_wire_834;
	wire [0 : 0] fresh_wire_835;
	wire [0 : 0] fresh_wire_836;
	wire [0 : 0] fresh_wire_837;
	wire [0 : 0] fresh_wire_838;
	wire [0 : 0] fresh_wire_839;
	wire [0 : 0] fresh_wire_840;
	wire [0 : 0] fresh_wire_841;
	wire [0 : 0] fresh_wire_842;
	wire [0 : 0] fresh_wire_843;
	wire [0 : 0] fresh_wire_844;
	wire [0 : 0] fresh_wire_845;
	wire [0 : 0] fresh_wire_846;
	wire [0 : 0] fresh_wire_847;
	wire [0 : 0] fresh_wire_848;
	wire [0 : 0] fresh_wire_849;
	wire [0 : 0] fresh_wire_850;
	wire [0 : 0] fresh_wire_851;
	wire [0 : 0] fresh_wire_852;
	wire [0 : 0] fresh_wire_853;
	wire [0 : 0] fresh_wire_854;
	wire [0 : 0] fresh_wire_855;
	wire [0 : 0] fresh_wire_856;
	wire [1 : 0] fresh_wire_857;
	wire [1 : 0] fresh_wire_858;
	wire [0 : 0] fresh_wire_859;
	wire [0 : 0] fresh_wire_860;
	wire [47 : 0] fresh_wire_861;
	wire [47 : 0] fresh_wire_862;
	wire [0 : 0] fresh_wire_863;
	wire [15 : 0] fresh_wire_864;
	wire [15 : 0] fresh_wire_865;
	wire [15 : 0] fresh_wire_866;
	wire [0 : 0] fresh_wire_867;
	wire [15 : 0] fresh_wire_868;
	wire [15 : 0] fresh_wire_869;
	wire [15 : 0] fresh_wire_870;
	wire [0 : 0] fresh_wire_871;
	wire [15 : 0] fresh_wire_872;
	wire [15 : 0] fresh_wire_873;
	wire [15 : 0] fresh_wire_874;
	wire [0 : 0] fresh_wire_875;
	wire [15 : 0] fresh_wire_876;
	wire [15 : 0] fresh_wire_877;
	wire [15 : 0] fresh_wire_878;
	wire [0 : 0] fresh_wire_879;
	wire [0 : 0] fresh_wire_880;
	wire [0 : 0] fresh_wire_881;
	wire [0 : 0] fresh_wire_882;
	wire [0 : 0] fresh_wire_883;
	wire [0 : 0] fresh_wire_884;
	wire [0 : 0] fresh_wire_885;
	wire [0 : 0] fresh_wire_886;
	wire [0 : 0] fresh_wire_887;
	wire [0 : 0] fresh_wire_888;
	wire [0 : 0] fresh_wire_889;
	wire [0 : 0] fresh_wire_890;
	wire [0 : 0] fresh_wire_891;
	wire [0 : 0] fresh_wire_892;
	wire [0 : 0] fresh_wire_893;
	wire [0 : 0] fresh_wire_894;
	wire [0 : 0] fresh_wire_895;
	wire [1 : 0] fresh_wire_896;
	wire [1 : 0] fresh_wire_897;
	wire [1 : 0] fresh_wire_898;
	wire [0 : 0] fresh_wire_899;
	wire [1 : 0] fresh_wire_900;
	wire [1 : 0] fresh_wire_901;
	wire [1 : 0] fresh_wire_902;
	wire [0 : 0] fresh_wire_903;
	wire [1 : 0] fresh_wire_904;
	wire [1 : 0] fresh_wire_905;
	wire [1 : 0] fresh_wire_906;
	wire [0 : 0] fresh_wire_907;
	wire [1 : 0] fresh_wire_908;
	wire [1 : 0] fresh_wire_909;
	wire [1 : 0] fresh_wire_910;
	wire [0 : 0] fresh_wire_911;
	wire [1 : 0] fresh_wire_912;
	wire [1 : 0] fresh_wire_913;
	wire [1 : 0] fresh_wire_914;
	wire [0 : 0] fresh_wire_915;
	wire [47 : 0] fresh_wire_916;
	wire [47 : 0] fresh_wire_917;
	wire [47 : 0] fresh_wire_918;
	wire [0 : 0] fresh_wire_919;
	wire [47 : 0] fresh_wire_920;
	wire [47 : 0] fresh_wire_921;
	wire [47 : 0] fresh_wire_922;
	wire [0 : 0] fresh_wire_923;
	wire [1 : 0] fresh_wire_924;
	wire [1 : 0] fresh_wire_925;
	wire [1 : 0] fresh_wire_926;
	wire [0 : 0] fresh_wire_927;
	wire [0 : 0] fresh_wire_928;
	wire [0 : 0] fresh_wire_929;
	wire [0 : 0] fresh_wire_930;
	wire [0 : 0] fresh_wire_931;
	wire [0 : 0] fresh_wire_932;
	wire [0 : 0] fresh_wire_933;
	wire [0 : 0] fresh_wire_934;
	wire [0 : 0] fresh_wire_935;
	wire [0 : 0] fresh_wire_936;
	wire [0 : 0] fresh_wire_937;
	wire [15 : 0] fresh_wire_938;
	wire [15 : 0] fresh_wire_939;
	wire [0 : 0] fresh_wire_940;
	wire [15 : 0] fresh_wire_941;
	wire [15 : 0] fresh_wire_942;
	wire [15 : 0] fresh_wire_943;
	wire [0 : 0] fresh_wire_944;
	wire [15 : 0] fresh_wire_945;
	wire [15 : 0] fresh_wire_946;
	wire [15 : 0] fresh_wire_947;
	wire [0 : 0] fresh_wire_948;
	wire [0 : 0] fresh_wire_949;
	wire [15 : 0] fresh_wire_950;
	wire [15 : 0] fresh_wire_951;
	wire [15 : 0] fresh_wire_952;
	wire [0 : 0] fresh_wire_953;
	wire [15 : 0] fresh_wire_954;
	wire [15 : 0] fresh_wire_955;
	wire [15 : 0] fresh_wire_956;
	wire [0 : 0] fresh_wire_957;
	wire [0 : 0] fresh_wire_958;
	wire [0 : 0] fresh_wire_959;
	wire [0 : 0] fresh_wire_960;
	wire [0 : 0] fresh_wire_961;
	wire [0 : 0] fresh_wire_962;
	wire [0 : 0] fresh_wire_963;
	wire [0 : 0] fresh_wire_964;
	wire [0 : 0] fresh_wire_965;
	wire [0 : 0] fresh_wire_966;
	wire [0 : 0] fresh_wire_967;
	wire [0 : 0] fresh_wire_968;
	wire [0 : 0] fresh_wire_969;
	wire [0 : 0] fresh_wire_970;
	wire [0 : 0] fresh_wire_971;
	wire [0 : 0] fresh_wire_972;
	wire [0 : 0] fresh_wire_973;
	wire [15 : 0] fresh_wire_974;
	wire [15 : 0] fresh_wire_975;
	wire [15 : 0] fresh_wire_976;
	wire [0 : 0] fresh_wire_977;
	wire [0 : 0] fresh_wire_978;
	wire [0 : 0] fresh_wire_979;
	wire [0 : 0] fresh_wire_980;
	wire [0 : 0] fresh_wire_981;
	wire [0 : 0] fresh_wire_982;
	wire [0 : 0] fresh_wire_983;
	wire [0 : 0] fresh_wire_984;
	wire [0 : 0] fresh_wire_985;
	wire [0 : 0] fresh_wire_986;
	wire [0 : 0] fresh_wire_987;
	wire [0 : 0] fresh_wire_988;
	wire [0 : 0] fresh_wire_989;
	wire [0 : 0] fresh_wire_990;
	wire [0 : 0] fresh_wire_991;
	wire [0 : 0] fresh_wire_992;
	wire [0 : 0] fresh_wire_993;
	wire [8 : 0] fresh_wire_994;
	wire [8 : 0] fresh_wire_995;
	wire [8 : 0] fresh_wire_996;
	wire [0 : 0] fresh_wire_997;
	wire [0 : 0] fresh_wire_998;
	wire [0 : 0] fresh_wire_999;
	wire [0 : 0] fresh_wire_1000;
	wire [0 : 0] fresh_wire_1001;
	wire [0 : 0] fresh_wire_1002;
	wire [0 : 0] fresh_wire_1003;
	wire [0 : 0] fresh_wire_1004;
	wire [0 : 0] fresh_wire_1005;
	wire [0 : 0] fresh_wire_1006;
	wire [8 : 0] fresh_wire_1007;
	wire [8 : 0] fresh_wire_1008;
	wire [8 : 0] fresh_wire_1009;
	wire [0 : 0] fresh_wire_1010;
	wire [0 : 0] fresh_wire_1011;
	wire [0 : 0] fresh_wire_1012;
	wire [0 : 0] fresh_wire_1013;
	wire [0 : 0] fresh_wire_1014;
	wire [0 : 0] fresh_wire_1015;
	wire [0 : 0] fresh_wire_1016;
	wire [0 : 0] fresh_wire_1017;
	wire [0 : 0] fresh_wire_1018;
	wire [0 : 0] fresh_wire_1019;
	wire [0 : 0] fresh_wire_1020;
	wire [8 : 0] fresh_wire_1021;
	wire [15 : 0] fresh_wire_1022;
	wire [8 : 0] fresh_wire_1023;
	wire [15 : 0] fresh_wire_1024;
	wire [0 : 0] fresh_wire_1025;
	wire [0 : 0] fresh_wire_1026;
	wire [0 : 0] fresh_wire_1027;
	wire [0 : 0] fresh_wire_1028;
	wire [0 : 0] fresh_wire_1029;
	wire [0 : 0] fresh_wire_1030;
	wire [0 : 0] fresh_wire_1031;
	wire [0 : 0] fresh_wire_1032;
	wire [0 : 0] fresh_wire_1033;
	wire [0 : 0] fresh_wire_1034;
	wire [0 : 0] fresh_wire_1035;
	wire [15 : 0] fresh_wire_1036;
	wire [15 : 0] fresh_wire_1037;
	wire [0 : 0] fresh_wire_1038;
	wire [15 : 0] fresh_wire_1039;
	wire [15 : 0] fresh_wire_1040;
	wire [15 : 0] fresh_wire_1041;
	wire [0 : 0] fresh_wire_1042;
	wire [15 : 0] fresh_wire_1043;
	wire [15 : 0] fresh_wire_1044;
	wire [15 : 0] fresh_wire_1045;
	wire [0 : 0] fresh_wire_1046;
	wire [0 : 0] fresh_wire_1047;
	wire [15 : 0] fresh_wire_1048;
	wire [15 : 0] fresh_wire_1049;
	wire [15 : 0] fresh_wire_1050;
	wire [0 : 0] fresh_wire_1051;
	wire [15 : 0] fresh_wire_1052;
	wire [15 : 0] fresh_wire_1053;
	wire [15 : 0] fresh_wire_1054;
	wire [0 : 0] fresh_wire_1055;
	wire [0 : 0] fresh_wire_1056;
	wire [0 : 0] fresh_wire_1057;
	wire [0 : 0] fresh_wire_1058;
	wire [0 : 0] fresh_wire_1059;
	wire [0 : 0] fresh_wire_1060;
	wire [0 : 0] fresh_wire_1061;
	wire [0 : 0] fresh_wire_1062;
	wire [0 : 0] fresh_wire_1063;
	wire [0 : 0] fresh_wire_1064;
	wire [0 : 0] fresh_wire_1065;
	wire [0 : 0] fresh_wire_1066;
	wire [0 : 0] fresh_wire_1067;
	wire [0 : 0] fresh_wire_1068;
	wire [0 : 0] fresh_wire_1069;
	wire [0 : 0] fresh_wire_1070;
	wire [0 : 0] fresh_wire_1071;
	wire [15 : 0] fresh_wire_1072;
	wire [15 : 0] fresh_wire_1073;
	wire [15 : 0] fresh_wire_1074;
	wire [0 : 0] fresh_wire_1075;
	wire [0 : 0] fresh_wire_1076;
	wire [0 : 0] fresh_wire_1077;
	wire [0 : 0] fresh_wire_1078;
	wire [0 : 0] fresh_wire_1079;
	wire [0 : 0] fresh_wire_1080;
	wire [0 : 0] fresh_wire_1081;
	wire [0 : 0] fresh_wire_1082;
	wire [0 : 0] fresh_wire_1083;
	wire [0 : 0] fresh_wire_1084;
	wire [0 : 0] fresh_wire_1085;
	wire [0 : 0] fresh_wire_1086;
	wire [0 : 0] fresh_wire_1087;
	wire [0 : 0] fresh_wire_1088;
	wire [0 : 0] fresh_wire_1089;
	wire [0 : 0] fresh_wire_1090;
	wire [0 : 0] fresh_wire_1091;
	wire [8 : 0] fresh_wire_1092;
	wire [8 : 0] fresh_wire_1093;
	wire [8 : 0] fresh_wire_1094;
	wire [0 : 0] fresh_wire_1095;
	wire [0 : 0] fresh_wire_1096;
	wire [0 : 0] fresh_wire_1097;
	wire [0 : 0] fresh_wire_1098;
	wire [0 : 0] fresh_wire_1099;
	wire [0 : 0] fresh_wire_1100;
	wire [0 : 0] fresh_wire_1101;
	wire [0 : 0] fresh_wire_1102;
	wire [0 : 0] fresh_wire_1103;
	wire [0 : 0] fresh_wire_1104;
	wire [8 : 0] fresh_wire_1105;
	wire [8 : 0] fresh_wire_1106;
	wire [8 : 0] fresh_wire_1107;
	wire [0 : 0] fresh_wire_1108;
	wire [0 : 0] fresh_wire_1109;
	wire [0 : 0] fresh_wire_1110;
	wire [0 : 0] fresh_wire_1111;
	wire [0 : 0] fresh_wire_1112;
	wire [0 : 0] fresh_wire_1113;
	wire [0 : 0] fresh_wire_1114;
	wire [0 : 0] fresh_wire_1115;
	wire [0 : 0] fresh_wire_1116;
	wire [0 : 0] fresh_wire_1117;
	wire [0 : 0] fresh_wire_1118;
	wire [8 : 0] fresh_wire_1119;
	wire [15 : 0] fresh_wire_1120;
	wire [8 : 0] fresh_wire_1121;
	wire [15 : 0] fresh_wire_1122;
	wire [0 : 0] fresh_wire_1123;
	wire [15 : 0] fresh_wire_1124;
	wire [15 : 0] fresh_wire_1125;
	wire [0 : 0] fresh_wire_1126;
	wire [0 : 0] fresh_wire_1127;
	wire [0 : 0] fresh_wire_1128;
	wire [0 : 0] fresh_wire_1129;
	wire [0 : 0] fresh_wire_1130;
	wire [0 : 0] fresh_wire_1131;
	wire [0 : 0] fresh_wire_1132;
	wire [0 : 0] fresh_wire_1133;
	wire [0 : 0] fresh_wire_1134;
	wire [0 : 0] fresh_wire_1135;
	wire [15 : 0] fresh_wire_1136;
	wire [15 : 0] fresh_wire_1137;
	wire [15 : 0] fresh_wire_1138;
	wire [1 : 0] fresh_wire_1139;
	wire [15 : 0] fresh_wire_1140;
	wire [15 : 0] fresh_wire_1141;
	wire [15 : 0] fresh_wire_1142;
	wire [15 : 0] fresh_wire_1143;
	wire [15 : 0] fresh_wire_1144;
	wire [31 : 0] fresh_wire_1145;
	wire [31 : 0] fresh_wire_1146;
	wire [31 : 0] fresh_wire_1147;
	wire [31 : 0] fresh_wire_1148;
	wire [15 : 0] fresh_wire_1149;
	wire [31 : 0] fresh_wire_1150;
	wire [31 : 0] fresh_wire_1151;
	wire [31 : 0] fresh_wire_1152;
	wire [31 : 0] fresh_wire_1153;
	wire [15 : 0] fresh_wire_1154;
	wire [31 : 0] fresh_wire_1155;
	wire [31 : 0] fresh_wire_1156;
	wire [31 : 0] fresh_wire_1157;
	wire [31 : 0] fresh_wire_1158;
	wire [15 : 0] fresh_wire_1159;
	wire [15 : 0] fresh_wire_1160;
	wire [15 : 0] fresh_wire_1161;
	wire [15 : 0] fresh_wire_1162;
	wire [15 : 0] fresh_wire_1163;
	wire [15 : 0] fresh_wire_1164;
	wire [15 : 0] fresh_wire_1165;
	wire [15 : 0] fresh_wire_1166;
	wire [15 : 0] fresh_wire_1167;
	wire [15 : 0] fresh_wire_1168;
	wire [15 : 0] fresh_wire_1169;
	wire [15 : 0] fresh_wire_1170;
	wire [0 : 0] fresh_wire_1171;
	wire [0 : 0] fresh_wire_1172;
	wire [0 : 0] fresh_wire_1173;
	wire [1 : 0] fresh_wire_1174;
	wire [1 : 0] fresh_wire_1175;
	wire [0 : 0] fresh_wire_1176;
	wire [1 : 0] fresh_wire_1177;
	wire [1 : 0] fresh_wire_1178;
	wire [0 : 0] fresh_wire_1179;
	wire [1 : 0] fresh_wire_1180;
	wire [1 : 0] fresh_wire_1181;
	wire [0 : 0] fresh_wire_1182;
	wire [15 : 0] fresh_wire_1183;
	wire [15 : 0] fresh_wire_1184;
	wire [0 : 0] fresh_wire_1185;
	wire [0 : 0] fresh_wire_1186;
	wire [0 : 0] fresh_wire_1187;
	wire [0 : 0] fresh_wire_1188;
	wire [0 : 0] fresh_wire_1189;
	wire [0 : 0] fresh_wire_1190;
	wire [0 : 0] fresh_wire_1191;
	wire [0 : 0] fresh_wire_1192;
	wire [0 : 0] fresh_wire_1193;
	wire [0 : 0] fresh_wire_1194;
	wire [0 : 0] fresh_wire_1195;
	wire [0 : 0] fresh_wire_1196;
	wire [0 : 0] fresh_wire_1197;
	wire [1 : 0] fresh_wire_1198;
	wire [1 : 0] fresh_wire_1199;
	wire [0 : 0] fresh_wire_1200;
	wire [0 : 0] fresh_wire_1201;
	wire [0 : 0] fresh_wire_1202;
	wire [0 : 0] fresh_wire_1203;
	wire [0 : 0] fresh_wire_1204;
	wire [0 : 0] fresh_wire_1205;
	wire [0 : 0] fresh_wire_1206;
	wire [1 : 0] fresh_wire_1207;
	wire [1 : 0] fresh_wire_1208;
	wire [0 : 0] fresh_wire_1209;
	wire [0 : 0] fresh_wire_1210;
	wire [0 : 0] fresh_wire_1211;
	wire [0 : 0] fresh_wire_1212;
	wire [0 : 0] fresh_wire_1213;
	wire [0 : 0] fresh_wire_1214;
	wire [0 : 0] fresh_wire_1215;
	wire [1 : 0] fresh_wire_1216;
	wire [1 : 0] fresh_wire_1217;
	wire [0 : 0] fresh_wire_1218;
	wire [1 : 0] fresh_wire_1219;
	wire [1 : 0] fresh_wire_1220;
	wire [0 : 0] fresh_wire_1221;
	wire [15 : 0] fresh_wire_1222;
	wire [15 : 0] fresh_wire_1223;
	wire [0 : 0] fresh_wire_1224;
	wire [0 : 0] fresh_wire_1225;
	wire [0 : 0] fresh_wire_1226;
	wire [0 : 0] fresh_wire_1227;
	wire [0 : 0] fresh_wire_1228;
	wire [0 : 0] fresh_wire_1229;
	wire [0 : 0] fresh_wire_1230;
	wire [15 : 0] fresh_wire_1231;
	wire [15 : 0] fresh_wire_1232;
	wire [0 : 0] fresh_wire_1233;
	wire [15 : 0] fresh_wire_1234;
	wire [15 : 0] fresh_wire_1235;
	wire [0 : 0] fresh_wire_1236;
	wire [15 : 0] fresh_wire_1237;
	wire [15 : 0] fresh_wire_1238;
	wire [0 : 0] fresh_wire_1239;
	wire [0 : 0] fresh_wire_1240;
	wire [0 : 0] fresh_wire_1241;
	wire [0 : 0] fresh_wire_1242;
	wire [0 : 0] fresh_wire_1243;
	wire [0 : 0] fresh_wire_1244;
	wire [0 : 0] fresh_wire_1245;
	wire [0 : 0] fresh_wire_1246;
	wire [0 : 0] fresh_wire_1247;
	wire [0 : 0] fresh_wire_1248;
	wire [0 : 0] fresh_wire_1249;
	wire [0 : 0] fresh_wire_1250;
	wire [0 : 0] fresh_wire_1251;
	wire [0 : 0] fresh_wire_1252;
	wire [0 : 0] fresh_wire_1253;
	wire [0 : 0] fresh_wire_1254;
	wire [0 : 0] fresh_wire_1255;
	wire [0 : 0] fresh_wire_1256;
	wire [0 : 0] fresh_wire_1257;
	wire [0 : 0] fresh_wire_1258;
	wire [0 : 0] fresh_wire_1259;
	wire [0 : 0] fresh_wire_1260;
	wire [0 : 0] fresh_wire_1261;
	wire [0 : 0] fresh_wire_1262;
	wire [0 : 0] fresh_wire_1263;
	wire [0 : 0] fresh_wire_1264;
	wire [0 : 0] fresh_wire_1265;
	wire [0 : 0] fresh_wire_1266;
	wire [0 : 0] fresh_wire_1267;
	wire [0 : 0] fresh_wire_1268;
	wire [0 : 0] fresh_wire_1269;
	wire [0 : 0] fresh_wire_1270;
	wire [0 : 0] fresh_wire_1271;
	wire [0 : 0] fresh_wire_1272;
	wire [0 : 0] fresh_wire_1273;
	wire [0 : 0] fresh_wire_1274;
	wire [0 : 0] fresh_wire_1275;
	wire [0 : 0] fresh_wire_1276;
	wire [0 : 0] fresh_wire_1277;
	wire [0 : 0] fresh_wire_1278;
	wire [0 : 0] fresh_wire_1279;
	wire [0 : 0] fresh_wire_1280;
	wire [0 : 0] fresh_wire_1281;
	wire [0 : 0] fresh_wire_1282;
	wire [0 : 0] fresh_wire_1283;
	wire [0 : 0] fresh_wire_1284;
	wire [0 : 0] fresh_wire_1285;
	wire [0 : 0] fresh_wire_1286;
	wire [0 : 0] fresh_wire_1287;
	wire [0 : 0] fresh_wire_1288;
	wire [0 : 0] fresh_wire_1289;
	wire [0 : 0] fresh_wire_1290;
	wire [0 : 0] fresh_wire_1291;
	wire [0 : 0] fresh_wire_1292;
	wire [0 : 0] fresh_wire_1293;
	wire [0 : 0] fresh_wire_1294;
	wire [0 : 0] fresh_wire_1295;
	wire [0 : 0] fresh_wire_1296;
	wire [0 : 0] fresh_wire_1297;
	wire [0 : 0] fresh_wire_1298;
	wire [0 : 0] fresh_wire_1299;
	wire [0 : 0] fresh_wire_1300;
	wire [0 : 0] fresh_wire_1301;
	wire [0 : 0] fresh_wire_1302;
	wire [0 : 0] fresh_wire_1303;
	wire [0 : 0] fresh_wire_1304;
	wire [0 : 0] fresh_wire_1305;
	wire [0 : 0] fresh_wire_1306;
	wire [0 : 0] fresh_wire_1307;
	wire [0 : 0] fresh_wire_1308;
	wire [0 : 0] fresh_wire_1309;
	wire [0 : 0] fresh_wire_1310;
	wire [0 : 0] fresh_wire_1311;
	wire [0 : 0] fresh_wire_1312;
	wire [0 : 0] fresh_wire_1313;
	wire [0 : 0] fresh_wire_1314;
	wire [0 : 0] fresh_wire_1315;
	wire [0 : 0] fresh_wire_1316;
	wire [0 : 0] fresh_wire_1317;
	wire [0 : 0] fresh_wire_1318;
	wire [0 : 0] fresh_wire_1319;
	wire [0 : 0] fresh_wire_1320;
	wire [0 : 0] fresh_wire_1321;
	wire [0 : 0] fresh_wire_1322;
	wire [0 : 0] fresh_wire_1323;
	wire [0 : 0] fresh_wire_1324;
	wire [0 : 0] fresh_wire_1325;
	wire [0 : 0] fresh_wire_1326;
	wire [0 : 0] fresh_wire_1327;
	wire [0 : 0] fresh_wire_1328;
	wire [0 : 0] fresh_wire_1329;
	wire [0 : 0] fresh_wire_1330;
	wire [0 : 0] fresh_wire_1331;
	wire [0 : 0] fresh_wire_1332;
	wire [15 : 0] fresh_wire_1333;
	wire [15 : 0] fresh_wire_1334;
	wire [0 : 0] fresh_wire_1335;
	wire [15 : 0] fresh_wire_1336;
	wire [15 : 0] fresh_wire_1337;
	wire [0 : 0] fresh_wire_1338;
	wire [0 : 0] fresh_wire_1339;
	wire [0 : 0] fresh_wire_1340;
	wire [0 : 0] fresh_wire_1341;
	wire [0 : 0] fresh_wire_1342;
	wire [0 : 0] fresh_wire_1343;
	wire [1 : 0] fresh_wire_1344;
	wire [1 : 0] fresh_wire_1345;
	wire [0 : 0] fresh_wire_1346;
	wire [1 : 0] fresh_wire_1347;
	wire [1 : 0] fresh_wire_1348;
	wire [0 : 0] fresh_wire_1349;
	wire [15 : 0] fresh_wire_1350;
	wire [15 : 0] fresh_wire_1351;
	wire [0 : 0] fresh_wire_1352;
	wire [0 : 0] fresh_wire_1353;
	wire [0 : 0] fresh_wire_1354;
	wire [0 : 0] fresh_wire_1355;
	wire [0 : 0] fresh_wire_1356;
	wire [0 : 0] fresh_wire_1357;
	wire [0 : 0] fresh_wire_1358;
	wire [0 : 0] fresh_wire_1359;
	wire [0 : 0] fresh_wire_1360;
	wire [0 : 0] fresh_wire_1361;
	wire [0 : 0] fresh_wire_1362;
	wire [0 : 0] fresh_wire_1363;
	wire [0 : 0] fresh_wire_1364;
	wire [0 : 0] fresh_wire_1365;
	wire [0 : 0] fresh_wire_1366;
	wire [0 : 0] fresh_wire_1367;
	wire [0 : 0] fresh_wire_1368;
	wire [0 : 0] fresh_wire_1369;
	wire [0 : 0] fresh_wire_1370;
	wire [0 : 0] fresh_wire_1371;
	wire [0 : 0] fresh_wire_1372;
	wire [1 : 0] fresh_wire_1373;
	wire [1 : 0] fresh_wire_1374;
	wire [0 : 0] fresh_wire_1375;
	wire [0 : 0] fresh_wire_1376;
	wire [15 : 0] fresh_wire_1377;
	wire [15 : 0] fresh_wire_1378;
	wire [0 : 0] fresh_wire_1379;
	wire [0 : 0] fresh_wire_1380;
	wire [15 : 0] fresh_wire_1381;
	wire [15 : 0] fresh_wire_1382;
	wire [0 : 0] fresh_wire_1383;
	wire [0 : 0] fresh_wire_1384;
	wire [15 : 0] fresh_wire_1385;
	wire [15 : 0] fresh_wire_1386;
	wire [0 : 0] fresh_wire_1387;
	wire [0 : 0] fresh_wire_1388;
	wire [15 : 0] fresh_wire_1389;
	wire [15 : 0] fresh_wire_1390;
	wire [0 : 0] fresh_wire_1391;
	wire [0 : 0] fresh_wire_1392;
	wire [0 : 0] fresh_wire_1393;
	wire [0 : 0] fresh_wire_1394;
	wire [0 : 0] fresh_wire_1395;
	wire [0 : 0] fresh_wire_1396;
	wire [0 : 0] fresh_wire_1397;
	wire [0 : 0] fresh_wire_1398;
	wire [0 : 0] fresh_wire_1399;
	wire [0 : 0] fresh_wire_1400;
	wire [0 : 0] fresh_wire_1401;
	wire [0 : 0] fresh_wire_1402;
	wire [0 : 0] fresh_wire_1403;
	wire [0 : 0] fresh_wire_1404;
	wire [15 : 0] fresh_wire_1405;
	wire [15 : 0] fresh_wire_1406;
	wire [15 : 0] fresh_wire_1407;
	wire [0 : 0] fresh_wire_1408;
	wire [0 : 0] fresh_wire_1409;
	wire [0 : 0] fresh_wire_1410;
	wire [0 : 0] fresh_wire_1411;
	wire [0 : 0] fresh_wire_1412;
	wire [0 : 0] fresh_wire_1413;
	wire [0 : 0] fresh_wire_1414;
	wire [0 : 0] fresh_wire_1415;
	wire [0 : 0] fresh_wire_1416;
	wire [0 : 0] fresh_wire_1417;
	wire [0 : 0] fresh_wire_1418;
	wire [0 : 0] fresh_wire_1419;
	wire [0 : 0] fresh_wire_1420;
	wire [0 : 0] fresh_wire_1421;
	wire [0 : 0] fresh_wire_1422;
	wire [0 : 0] fresh_wire_1423;
	wire [0 : 0] fresh_wire_1424;
	wire [0 : 0] fresh_wire_1425;
	wire [0 : 0] fresh_wire_1426;
	wire [0 : 0] fresh_wire_1427;
	wire [0 : 0] fresh_wire_1428;
	wire [15 : 0] fresh_wire_1429;
	wire [15 : 0] fresh_wire_1430;
	wire [15 : 0] fresh_wire_1431;
	wire [0 : 0] fresh_wire_1432;
	wire [15 : 0] fresh_wire_1433;
	wire [15 : 0] fresh_wire_1434;
	wire [15 : 0] fresh_wire_1435;
	wire [0 : 0] fresh_wire_1436;
	wire [15 : 0] fresh_wire_1437;
	wire [15 : 0] fresh_wire_1438;
	wire [15 : 0] fresh_wire_1439;
	wire [0 : 0] fresh_wire_1440;
	wire [15 : 0] fresh_wire_1441;
	wire [15 : 0] fresh_wire_1442;
	wire [15 : 0] fresh_wire_1443;
	wire [0 : 0] fresh_wire_1444;
	wire [1 : 0] fresh_wire_1445;
	wire [1 : 0] fresh_wire_1446;
	wire [1 : 0] fresh_wire_1447;
	wire [0 : 0] fresh_wire_1448;
	wire [1 : 0] fresh_wire_1449;
	wire [1 : 0] fresh_wire_1450;
	wire [1 : 0] fresh_wire_1451;
	wire [0 : 0] fresh_wire_1452;
	wire [1 : 0] fresh_wire_1453;
	wire [1 : 0] fresh_wire_1454;
	wire [1 : 0] fresh_wire_1455;
	wire [0 : 0] fresh_wire_1456;
	wire [1 : 0] fresh_wire_1457;
	wire [1 : 0] fresh_wire_1458;
	wire [1 : 0] fresh_wire_1459;
	wire [0 : 0] fresh_wire_1460;
	wire [1 : 0] fresh_wire_1461;
	wire [1 : 0] fresh_wire_1462;
	wire [1 : 0] fresh_wire_1463;
	wire [0 : 0] fresh_wire_1464;
	wire [1 : 0] fresh_wire_1465;
	wire [1 : 0] fresh_wire_1466;
	wire [1 : 0] fresh_wire_1467;
	wire [0 : 0] fresh_wire_1468;
	wire [0 : 0] fresh_wire_1469;
	wire [0 : 0] fresh_wire_1470;
	wire [0 : 0] fresh_wire_1471;
	wire [0 : 0] fresh_wire_1472;
	wire [0 : 0] fresh_wire_1473;
	wire [0 : 0] fresh_wire_1474;
	wire [0 : 0] fresh_wire_1475;
	wire [0 : 0] fresh_wire_1476;
	wire [0 : 0] fresh_wire_1477;
	wire [0 : 0] fresh_wire_1478;
	wire [0 : 0] fresh_wire_1479;
	wire [0 : 0] fresh_wire_1480;
	wire [0 : 0] fresh_wire_1481;
	wire [0 : 0] fresh_wire_1482;
	wire [0 : 0] fresh_wire_1483;
	wire [0 : 0] fresh_wire_1484;
	wire [0 : 0] fresh_wire_1485;
	wire [0 : 0] fresh_wire_1486;
	wire [0 : 0] fresh_wire_1487;
	wire [0 : 0] fresh_wire_1488;
	wire [0 : 0] fresh_wire_1489;
	wire [0 : 0] fresh_wire_1490;
	wire [0 : 0] fresh_wire_1491;
	wire [0 : 0] fresh_wire_1492;
	wire [0 : 0] fresh_wire_1493;
	wire [0 : 0] fresh_wire_1494;
	wire [0 : 0] fresh_wire_1495;
	wire [0 : 0] fresh_wire_1496;
	wire [0 : 0] fresh_wire_1497;
	wire [0 : 0] fresh_wire_1498;
	wire [0 : 0] fresh_wire_1499;
	wire [0 : 0] fresh_wire_1500;
	wire [0 : 0] fresh_wire_1501;
	wire [0 : 0] fresh_wire_1502;
	wire [0 : 0] fresh_wire_1503;
	wire [0 : 0] fresh_wire_1504;
	wire [0 : 0] fresh_wire_1505;
	wire [0 : 0] fresh_wire_1506;
	wire [0 : 0] fresh_wire_1507;
	wire [0 : 0] fresh_wire_1508;
	wire [15 : 0] fresh_wire_1509;
	wire [15 : 0] fresh_wire_1510;
	wire [15 : 0] fresh_wire_1511;
	wire [0 : 0] fresh_wire_1512;
	wire [15 : 0] fresh_wire_1513;
	wire [15 : 0] fresh_wire_1514;
	wire [15 : 0] fresh_wire_1515;
	wire [0 : 0] fresh_wire_1516;
	wire [15 : 0] fresh_wire_1517;
	wire [15 : 0] fresh_wire_1518;
	wire [15 : 0] fresh_wire_1519;
	wire [0 : 0] fresh_wire_1520;
	wire [15 : 0] fresh_wire_1521;
	wire [15 : 0] fresh_wire_1522;
	wire [15 : 0] fresh_wire_1523;
	wire [0 : 0] fresh_wire_1524;
	wire [15 : 0] fresh_wire_1525;
	wire [15 : 0] fresh_wire_1526;
	wire [15 : 0] fresh_wire_1527;
	wire [0 : 0] fresh_wire_1528;
	wire [15 : 0] fresh_wire_1529;
	wire [15 : 0] fresh_wire_1530;
	wire [15 : 0] fresh_wire_1531;
	wire [0 : 0] fresh_wire_1532;
	wire [15 : 0] fresh_wire_1533;
	wire [15 : 0] fresh_wire_1534;
	wire [15 : 0] fresh_wire_1535;
	wire [0 : 0] fresh_wire_1536;
	wire [15 : 0] fresh_wire_1537;
	wire [15 : 0] fresh_wire_1538;
	wire [15 : 0] fresh_wire_1539;
	wire [0 : 0] fresh_wire_1540;
	wire [15 : 0] fresh_wire_1541;
	wire [15 : 0] fresh_wire_1542;
	wire [15 : 0] fresh_wire_1543;
	wire [0 : 0] fresh_wire_1544;
	wire [0 : 0] fresh_wire_1545;
	wire [0 : 0] fresh_wire_1546;
	wire [0 : 0] fresh_wire_1547;
	wire [0 : 0] fresh_wire_1548;
	wire [0 : 0] fresh_wire_1549;
	wire [0 : 0] fresh_wire_1550;
	wire [0 : 0] fresh_wire_1551;
	wire [0 : 0] fresh_wire_1552;
	wire [0 : 0] fresh_wire_1553;
	wire [0 : 0] fresh_wire_1554;
	wire [0 : 0] fresh_wire_1555;
	wire [0 : 0] fresh_wire_1556;
	wire [0 : 0] fresh_wire_1557;
	wire [0 : 0] fresh_wire_1558;
	wire [0 : 0] fresh_wire_1559;
	wire [0 : 0] fresh_wire_1560;
	wire [0 : 0] fresh_wire_1561;
	wire [0 : 0] fresh_wire_1562;
	wire [0 : 0] fresh_wire_1563;
	wire [0 : 0] fresh_wire_1564;
	wire [15 : 0] fresh_wire_1565;
	wire [31 : 0] fresh_wire_1566;
	wire [31 : 0] fresh_wire_1567;
	wire [31 : 0] fresh_wire_1568;
	wire [31 : 0] fresh_wire_1569;
	wire [31 : 0] fresh_wire_1570;
	wire [31 : 0] fresh_wire_1571;
	wire [31 : 0] fresh_wire_1572;
	wire [0 : 0] fresh_wire_1573;
	wire [15 : 0] fresh_wire_1574;
	wire [15 : 0] fresh_wire_1575;
	wire [15 : 0] fresh_wire_1576;
	wire [0 : 0] fresh_wire_1577;
	wire [0 : 0] fresh_wire_1578;
	wire [15 : 0] fresh_wire_1579;
	wire [15 : 0] fresh_wire_1580;
	wire [15 : 0] fresh_wire_1581;
	wire [0 : 0] fresh_wire_1582;
	wire [1 : 0] fresh_wire_1583;
	wire [1 : 0] fresh_wire_1584;
	wire [1 : 0] fresh_wire_1585;
	wire [0 : 0] fresh_wire_1586;
	wire [0 : 0] fresh_wire_1587;
	wire [0 : 0] fresh_wire_1588;
	wire [0 : 0] fresh_wire_1589;
	wire [0 : 0] fresh_wire_1590;
	wire [0 : 0] fresh_wire_1591;
	wire [0 : 0] fresh_wire_1592;
	wire [0 : 0] fresh_wire_1593;
	wire [0 : 0] fresh_wire_1594;
	wire [1 : 0] fresh_wire_1595;
	wire [1 : 0] fresh_wire_1596;
	wire [0 : 0] fresh_wire_1597;
	wire [1 : 0] fresh_wire_1598;
	wire [1 : 0] fresh_wire_1599;
	wire [0 : 0] fresh_wire_1600;
	wire [0 : 0] fresh_wire_1601;
	wire [0 : 0] fresh_wire_1602;
	wire [0 : 0] fresh_wire_1603;
	wire [1 : 0] fresh_wire_1604;
	wire [1 : 0] fresh_wire_1605;
	wire [0 : 0] fresh_wire_1606;
	wire [1 : 0] fresh_wire_1607;
	wire [1 : 0] fresh_wire_1608;
	wire [0 : 0] fresh_wire_1609;
	wire [0 : 0] fresh_wire_1610;
	wire [0 : 0] fresh_wire_1611;
	wire [0 : 0] fresh_wire_1612;
	wire [0 : 0] fresh_wire_1613;
	wire [0 : 0] fresh_wire_1614;
	wire [0 : 0] fresh_wire_1615;
	wire [0 : 0] fresh_wire_1616;
	wire [0 : 0] fresh_wire_1617;
	wire [0 : 0] fresh_wire_1618;
	wire [0 : 0] fresh_wire_1619;
	wire [0 : 0] fresh_wire_1620;
	wire [0 : 0] fresh_wire_1621;
	wire [0 : 0] fresh_wire_1622;
	wire [0 : 0] fresh_wire_1623;
	wire [0 : 0] fresh_wire_1624;
	wire [0 : 0] fresh_wire_1625;
	wire [0 : 0] fresh_wire_1626;
	wire [0 : 0] fresh_wire_1627;
	wire [0 : 0] fresh_wire_1628;
	wire [0 : 0] fresh_wire_1629;
	wire [0 : 0] fresh_wire_1630;
	wire [0 : 0] fresh_wire_1631;
	wire [0 : 0] fresh_wire_1632;
	wire [0 : 0] fresh_wire_1633;
	wire [0 : 0] fresh_wire_1634;
	wire [0 : 0] fresh_wire_1635;
	wire [0 : 0] fresh_wire_1636;
	wire [1 : 0] fresh_wire_1637;
	wire [1 : 0] fresh_wire_1638;
	wire [0 : 0] fresh_wire_1639;
	wire [0 : 0] fresh_wire_1640;
	wire [47 : 0] fresh_wire_1641;
	wire [47 : 0] fresh_wire_1642;
	wire [0 : 0] fresh_wire_1643;
	wire [0 : 0] fresh_wire_1644;
	wire [0 : 0] fresh_wire_1645;
	wire [0 : 0] fresh_wire_1646;
	wire [0 : 0] fresh_wire_1647;
	wire [0 : 0] fresh_wire_1648;
	wire [0 : 0] fresh_wire_1649;
	wire [0 : 0] fresh_wire_1650;
	wire [0 : 0] fresh_wire_1651;
	wire [1 : 0] fresh_wire_1652;
	wire [1 : 0] fresh_wire_1653;
	wire [1 : 0] fresh_wire_1654;
	wire [0 : 0] fresh_wire_1655;
	wire [1 : 0] fresh_wire_1656;
	wire [1 : 0] fresh_wire_1657;
	wire [1 : 0] fresh_wire_1658;
	wire [0 : 0] fresh_wire_1659;
	wire [31 : 0] fresh_wire_1660;
	wire [31 : 0] fresh_wire_1661;
	wire [31 : 0] fresh_wire_1662;
	wire [0 : 0] fresh_wire_1663;
	wire [31 : 0] fresh_wire_1664;
	wire [31 : 0] fresh_wire_1665;
	wire [31 : 0] fresh_wire_1666;
	wire [0 : 0] fresh_wire_1667;
	wire [31 : 0] fresh_wire_1668;
	wire [31 : 0] fresh_wire_1669;
	wire [31 : 0] fresh_wire_1670;
	wire [0 : 0] fresh_wire_1671;
	wire [31 : 0] fresh_wire_1672;
	wire [31 : 0] fresh_wire_1673;
	wire [31 : 0] fresh_wire_1674;
	wire [0 : 0] fresh_wire_1675;
	wire [31 : 0] fresh_wire_1676;
	wire [31 : 0] fresh_wire_1677;
	wire [31 : 0] fresh_wire_1678;
	wire [0 : 0] fresh_wire_1679;
	wire [31 : 0] fresh_wire_1680;
	wire [31 : 0] fresh_wire_1681;
	wire [31 : 0] fresh_wire_1682;
	wire [0 : 0] fresh_wire_1683;
	wire [31 : 0] fresh_wire_1684;
	wire [31 : 0] fresh_wire_1685;
	wire [31 : 0] fresh_wire_1686;
	wire [0 : 0] fresh_wire_1687;
	wire [1 : 0] fresh_wire_1688;
	wire [1 : 0] fresh_wire_1689;
	wire [1 : 0] fresh_wire_1690;
	wire [0 : 0] fresh_wire_1691;
	wire [1 : 0] fresh_wire_1692;
	wire [1 : 0] fresh_wire_1693;
	wire [1 : 0] fresh_wire_1694;
	wire [1 : 0] fresh_wire_1695;
	wire [1 : 0] fresh_wire_1696;
	wire [1 : 0] fresh_wire_1697;
	wire [0 : 0] fresh_wire_1698;
	wire [0 : 0] fresh_wire_1699;
	wire [0 : 0] fresh_wire_1700;
	wire [0 : 0] fresh_wire_1701;
	wire [0 : 0] fresh_wire_1702;
	wire [0 : 0] fresh_wire_1703;
	wire [0 : 0] fresh_wire_1704;
	wire [0 : 0] fresh_wire_1705;
	wire [0 : 0] fresh_wire_1706;
	wire [0 : 0] fresh_wire_1707;
	wire [0 : 0] fresh_wire_1708;
	wire [0 : 0] fresh_wire_1709;
	wire [0 : 0] fresh_wire_1710;
	wire [0 : 0] fresh_wire_1711;
	wire [0 : 0] fresh_wire_1712;
	wire [0 : 0] fresh_wire_1713;
	wire [0 : 0] fresh_wire_1714;
	wire [0 : 0] fresh_wire_1715;
	wire [1 : 0] fresh_wire_1716;
	wire [1 : 0] fresh_wire_1717;
	wire [0 : 0] fresh_wire_1718;
	wire [1 : 0] fresh_wire_1719;
	wire [1 : 0] fresh_wire_1720;
	wire [0 : 0] fresh_wire_1721;
	wire [1 : 0] fresh_wire_1722;
	wire [1 : 0] fresh_wire_1723;
	wire [0 : 0] fresh_wire_1724;
	wire [1 : 0] fresh_wire_1725;
	wire [1 : 0] fresh_wire_1726;
	wire [0 : 0] fresh_wire_1727;
	wire [1 : 0] fresh_wire_1728;
	wire [1 : 0] fresh_wire_1729;
	wire [0 : 0] fresh_wire_1730;
	wire [0 : 0] fresh_wire_1731;
	wire [0 : 0] fresh_wire_1732;
	wire [0 : 0] fresh_wire_1733;
	wire [0 : 0] fresh_wire_1734;
	wire [0 : 0] fresh_wire_1735;
	wire [0 : 0] fresh_wire_1736;
	wire [0 : 0] fresh_wire_1737;
	wire [0 : 0] fresh_wire_1738;
	wire [0 : 0] fresh_wire_1739;
	wire [0 : 0] fresh_wire_1740;
	wire [0 : 0] fresh_wire_1741;
	wire [0 : 0] fresh_wire_1742;
	wire [0 : 0] fresh_wire_1743;
	wire [0 : 0] fresh_wire_1744;
	wire [0 : 0] fresh_wire_1745;
	wire [0 : 0] fresh_wire_1746;
	wire [0 : 0] fresh_wire_1747;
	wire [0 : 0] fresh_wire_1748;
	wire [0 : 0] fresh_wire_1749;
	wire [0 : 0] fresh_wire_1750;
	wire [0 : 0] fresh_wire_1751;
	wire [0 : 0] fresh_wire_1752;
	wire [0 : 0] fresh_wire_1753;
	wire [0 : 0] fresh_wire_1754;
	wire [0 : 0] fresh_wire_1755;
	wire [0 : 0] fresh_wire_1756;
	wire [0 : 0] fresh_wire_1757;
	wire [0 : 0] fresh_wire_1758;
	wire [0 : 0] fresh_wire_1759;
	wire [0 : 0] fresh_wire_1760;
	wire [0 : 0] fresh_wire_1761;
	wire [0 : 0] fresh_wire_1762;
	wire [0 : 0] fresh_wire_1763;
	wire [0 : 0] fresh_wire_1764;
	wire [0 : 0] fresh_wire_1765;
	wire [0 : 0] fresh_wire_1766;
	wire [0 : 0] fresh_wire_1767;
	wire [0 : 0] fresh_wire_1768;
	wire [0 : 0] fresh_wire_1769;
	wire [0 : 0] fresh_wire_1770;
	wire [0 : 0] fresh_wire_1771;
	wire [0 : 0] fresh_wire_1772;
	wire [0 : 0] fresh_wire_1773;
	wire [0 : 0] fresh_wire_1774;
	wire [0 : 0] fresh_wire_1775;
	wire [0 : 0] fresh_wire_1776;
	wire [0 : 0] fresh_wire_1777;
	wire [0 : 0] fresh_wire_1778;
	wire [0 : 0] fresh_wire_1779;
	wire [0 : 0] fresh_wire_1780;
	wire [0 : 0] fresh_wire_1781;
	wire [0 : 0] fresh_wire_1782;
	wire [0 : 0] fresh_wire_1783;
	wire [0 : 0] fresh_wire_1784;
	wire [0 : 0] fresh_wire_1785;
	wire [0 : 0] fresh_wire_1786;
	wire [0 : 0] fresh_wire_1787;
	wire [0 : 0] fresh_wire_1788;
	wire [0 : 0] fresh_wire_1789;
	wire [0 : 0] fresh_wire_1790;
	wire [0 : 0] fresh_wire_1791;
	wire [0 : 0] fresh_wire_1792;
	wire [0 : 0] fresh_wire_1793;
	wire [0 : 0] fresh_wire_1794;
	wire [0 : 0] fresh_wire_1795;
	wire [0 : 0] fresh_wire_1796;
	wire [0 : 0] fresh_wire_1797;
	wire [0 : 0] fresh_wire_1798;
	wire [0 : 0] fresh_wire_1799;
	wire [0 : 0] fresh_wire_1800;
	wire [0 : 0] fresh_wire_1801;
	wire [0 : 0] fresh_wire_1802;
	wire [0 : 0] fresh_wire_1803;
	wire [0 : 0] fresh_wire_1804;
	wire [0 : 0] fresh_wire_1805;
	wire [0 : 0] fresh_wire_1806;
	wire [0 : 0] fresh_wire_1807;
	wire [0 : 0] fresh_wire_1808;
	wire [0 : 0] fresh_wire_1809;
	wire [0 : 0] fresh_wire_1810;
	wire [0 : 0] fresh_wire_1811;
	wire [0 : 0] fresh_wire_1812;
	wire [0 : 0] fresh_wire_1813;
	wire [0 : 0] fresh_wire_1814;
	wire [0 : 0] fresh_wire_1815;
	wire [0 : 0] fresh_wire_1816;
	wire [0 : 0] fresh_wire_1817;
	wire [0 : 0] fresh_wire_1818;
	wire [0 : 0] fresh_wire_1819;
	wire [0 : 0] fresh_wire_1820;
	wire [0 : 0] fresh_wire_1821;
	wire [0 : 0] fresh_wire_1822;
	wire [0 : 0] fresh_wire_1823;
	wire [0 : 0] fresh_wire_1824;
	wire [0 : 0] fresh_wire_1825;
	wire [0 : 0] fresh_wire_1826;
	wire [0 : 0] fresh_wire_1827;
	wire [0 : 0] fresh_wire_1828;
	wire [1 : 0] fresh_wire_1829;
	wire [1 : 0] fresh_wire_1830;
	wire [0 : 0] fresh_wire_1831;
	wire [0 : 0] fresh_wire_1832;
	wire [47 : 0] fresh_wire_1833;
	wire [47 : 0] fresh_wire_1834;
	wire [0 : 0] fresh_wire_1835;
	wire [15 : 0] fresh_wire_1836;
	wire [15 : 0] fresh_wire_1837;
	wire [15 : 0] fresh_wire_1838;
	wire [0 : 0] fresh_wire_1839;
	wire [15 : 0] fresh_wire_1840;
	wire [15 : 0] fresh_wire_1841;
	wire [15 : 0] fresh_wire_1842;
	wire [0 : 0] fresh_wire_1843;
	wire [15 : 0] fresh_wire_1844;
	wire [15 : 0] fresh_wire_1845;
	wire [15 : 0] fresh_wire_1846;
	wire [0 : 0] fresh_wire_1847;
	wire [15 : 0] fresh_wire_1848;
	wire [15 : 0] fresh_wire_1849;
	wire [15 : 0] fresh_wire_1850;
	wire [0 : 0] fresh_wire_1851;
	wire [0 : 0] fresh_wire_1852;
	wire [0 : 0] fresh_wire_1853;
	wire [0 : 0] fresh_wire_1854;
	wire [0 : 0] fresh_wire_1855;
	wire [0 : 0] fresh_wire_1856;
	wire [0 : 0] fresh_wire_1857;
	wire [0 : 0] fresh_wire_1858;
	wire [0 : 0] fresh_wire_1859;
	wire [0 : 0] fresh_wire_1860;
	wire [0 : 0] fresh_wire_1861;
	wire [0 : 0] fresh_wire_1862;
	wire [0 : 0] fresh_wire_1863;
	wire [0 : 0] fresh_wire_1864;
	wire [0 : 0] fresh_wire_1865;
	wire [0 : 0] fresh_wire_1866;
	wire [0 : 0] fresh_wire_1867;
	wire [1 : 0] fresh_wire_1868;
	wire [1 : 0] fresh_wire_1869;
	wire [1 : 0] fresh_wire_1870;
	wire [0 : 0] fresh_wire_1871;
	wire [1 : 0] fresh_wire_1872;
	wire [1 : 0] fresh_wire_1873;
	wire [1 : 0] fresh_wire_1874;
	wire [0 : 0] fresh_wire_1875;
	wire [1 : 0] fresh_wire_1876;
	wire [1 : 0] fresh_wire_1877;
	wire [1 : 0] fresh_wire_1878;
	wire [0 : 0] fresh_wire_1879;
	wire [1 : 0] fresh_wire_1880;
	wire [1 : 0] fresh_wire_1881;
	wire [1 : 0] fresh_wire_1882;
	wire [0 : 0] fresh_wire_1883;
	wire [1 : 0] fresh_wire_1884;
	wire [1 : 0] fresh_wire_1885;
	wire [1 : 0] fresh_wire_1886;
	wire [0 : 0] fresh_wire_1887;
	wire [47 : 0] fresh_wire_1888;
	wire [47 : 0] fresh_wire_1889;
	wire [47 : 0] fresh_wire_1890;
	wire [0 : 0] fresh_wire_1891;
	wire [47 : 0] fresh_wire_1892;
	wire [47 : 0] fresh_wire_1893;
	wire [47 : 0] fresh_wire_1894;
	wire [0 : 0] fresh_wire_1895;
	wire [1 : 0] fresh_wire_1896;
	wire [1 : 0] fresh_wire_1897;
	wire [1 : 0] fresh_wire_1898;
	wire [0 : 0] fresh_wire_1899;
	wire [0 : 0] fresh_wire_1900;
	wire [0 : 0] fresh_wire_1901;
	wire [0 : 0] fresh_wire_1902;
	wire [0 : 0] fresh_wire_1903;
	wire [0 : 0] fresh_wire_1904;
	wire [0 : 0] fresh_wire_1905;
	wire [0 : 0] fresh_wire_1906;
	wire [0 : 0] fresh_wire_1907;
	wire [0 : 0] fresh_wire_1908;
	wire [0 : 0] fresh_wire_1909;
	wire [15 : 0] fresh_wire_1910;
	wire [15 : 0] fresh_wire_1911;
	wire [0 : 0] fresh_wire_1912;
	wire [15 : 0] fresh_wire_1913;
	wire [15 : 0] fresh_wire_1914;
	wire [15 : 0] fresh_wire_1915;
	wire [0 : 0] fresh_wire_1916;
	wire [15 : 0] fresh_wire_1917;
	wire [15 : 0] fresh_wire_1918;
	wire [15 : 0] fresh_wire_1919;
	wire [0 : 0] fresh_wire_1920;
	wire [0 : 0] fresh_wire_1921;
	wire [15 : 0] fresh_wire_1922;
	wire [15 : 0] fresh_wire_1923;
	wire [15 : 0] fresh_wire_1924;
	wire [0 : 0] fresh_wire_1925;
	wire [15 : 0] fresh_wire_1926;
	wire [15 : 0] fresh_wire_1927;
	wire [15 : 0] fresh_wire_1928;
	wire [0 : 0] fresh_wire_1929;
	wire [0 : 0] fresh_wire_1930;
	wire [0 : 0] fresh_wire_1931;
	wire [0 : 0] fresh_wire_1932;
	wire [0 : 0] fresh_wire_1933;
	wire [0 : 0] fresh_wire_1934;
	wire [0 : 0] fresh_wire_1935;
	wire [0 : 0] fresh_wire_1936;
	wire [0 : 0] fresh_wire_1937;
	wire [0 : 0] fresh_wire_1938;
	wire [0 : 0] fresh_wire_1939;
	wire [0 : 0] fresh_wire_1940;
	wire [0 : 0] fresh_wire_1941;
	wire [0 : 0] fresh_wire_1942;
	wire [0 : 0] fresh_wire_1943;
	wire [0 : 0] fresh_wire_1944;
	wire [0 : 0] fresh_wire_1945;
	wire [15 : 0] fresh_wire_1946;
	wire [15 : 0] fresh_wire_1947;
	wire [15 : 0] fresh_wire_1948;
	wire [0 : 0] fresh_wire_1949;
	wire [0 : 0] fresh_wire_1950;
	wire [0 : 0] fresh_wire_1951;
	wire [0 : 0] fresh_wire_1952;
	wire [0 : 0] fresh_wire_1953;
	wire [0 : 0] fresh_wire_1954;
	wire [0 : 0] fresh_wire_1955;
	wire [0 : 0] fresh_wire_1956;
	wire [0 : 0] fresh_wire_1957;
	wire [0 : 0] fresh_wire_1958;
	wire [0 : 0] fresh_wire_1959;
	wire [0 : 0] fresh_wire_1960;
	wire [0 : 0] fresh_wire_1961;
	wire [0 : 0] fresh_wire_1962;
	wire [0 : 0] fresh_wire_1963;
	wire [0 : 0] fresh_wire_1964;
	wire [0 : 0] fresh_wire_1965;
	wire [8 : 0] fresh_wire_1966;
	wire [8 : 0] fresh_wire_1967;
	wire [8 : 0] fresh_wire_1968;
	wire [0 : 0] fresh_wire_1969;
	wire [0 : 0] fresh_wire_1970;
	wire [0 : 0] fresh_wire_1971;
	wire [0 : 0] fresh_wire_1972;
	wire [0 : 0] fresh_wire_1973;
	wire [0 : 0] fresh_wire_1974;
	wire [0 : 0] fresh_wire_1975;
	wire [0 : 0] fresh_wire_1976;
	wire [0 : 0] fresh_wire_1977;
	wire [0 : 0] fresh_wire_1978;
	wire [8 : 0] fresh_wire_1979;
	wire [8 : 0] fresh_wire_1980;
	wire [8 : 0] fresh_wire_1981;
	wire [0 : 0] fresh_wire_1982;
	wire [0 : 0] fresh_wire_1983;
	wire [0 : 0] fresh_wire_1984;
	wire [0 : 0] fresh_wire_1985;
	wire [0 : 0] fresh_wire_1986;
	wire [0 : 0] fresh_wire_1987;
	wire [0 : 0] fresh_wire_1988;
	wire [0 : 0] fresh_wire_1989;
	wire [0 : 0] fresh_wire_1990;
	wire [0 : 0] fresh_wire_1991;
	wire [0 : 0] fresh_wire_1992;
	wire [8 : 0] fresh_wire_1993;
	wire [15 : 0] fresh_wire_1994;
	wire [8 : 0] fresh_wire_1995;
	wire [15 : 0] fresh_wire_1996;
	wire [0 : 0] fresh_wire_1997;
	wire [0 : 0] fresh_wire_1998;
	wire [0 : 0] fresh_wire_1999;
	wire [0 : 0] fresh_wire_2000;
	wire [0 : 0] fresh_wire_2001;
	wire [0 : 0] fresh_wire_2002;
	wire [0 : 0] fresh_wire_2003;
	wire [0 : 0] fresh_wire_2004;
	wire [0 : 0] fresh_wire_2005;
	wire [0 : 0] fresh_wire_2006;
	wire [0 : 0] fresh_wire_2007;
	wire [15 : 0] fresh_wire_2008;
	wire [15 : 0] fresh_wire_2009;
	wire [0 : 0] fresh_wire_2010;
	wire [15 : 0] fresh_wire_2011;
	wire [15 : 0] fresh_wire_2012;
	wire [15 : 0] fresh_wire_2013;
	wire [0 : 0] fresh_wire_2014;
	wire [15 : 0] fresh_wire_2015;
	wire [15 : 0] fresh_wire_2016;
	wire [15 : 0] fresh_wire_2017;
	wire [0 : 0] fresh_wire_2018;
	wire [0 : 0] fresh_wire_2019;
	wire [15 : 0] fresh_wire_2020;
	wire [15 : 0] fresh_wire_2021;
	wire [15 : 0] fresh_wire_2022;
	wire [0 : 0] fresh_wire_2023;
	wire [15 : 0] fresh_wire_2024;
	wire [15 : 0] fresh_wire_2025;
	wire [15 : 0] fresh_wire_2026;
	wire [0 : 0] fresh_wire_2027;
	wire [0 : 0] fresh_wire_2028;
	wire [0 : 0] fresh_wire_2029;
	wire [0 : 0] fresh_wire_2030;
	wire [0 : 0] fresh_wire_2031;
	wire [0 : 0] fresh_wire_2032;
	wire [0 : 0] fresh_wire_2033;
	wire [0 : 0] fresh_wire_2034;
	wire [0 : 0] fresh_wire_2035;
	wire [0 : 0] fresh_wire_2036;
	wire [0 : 0] fresh_wire_2037;
	wire [0 : 0] fresh_wire_2038;
	wire [0 : 0] fresh_wire_2039;
	wire [0 : 0] fresh_wire_2040;
	wire [0 : 0] fresh_wire_2041;
	wire [0 : 0] fresh_wire_2042;
	wire [0 : 0] fresh_wire_2043;
	wire [15 : 0] fresh_wire_2044;
	wire [15 : 0] fresh_wire_2045;
	wire [15 : 0] fresh_wire_2046;
	wire [0 : 0] fresh_wire_2047;
	wire [0 : 0] fresh_wire_2048;
	wire [0 : 0] fresh_wire_2049;
	wire [0 : 0] fresh_wire_2050;
	wire [0 : 0] fresh_wire_2051;
	wire [0 : 0] fresh_wire_2052;
	wire [0 : 0] fresh_wire_2053;
	wire [0 : 0] fresh_wire_2054;
	wire [0 : 0] fresh_wire_2055;
	wire [0 : 0] fresh_wire_2056;
	wire [0 : 0] fresh_wire_2057;
	wire [0 : 0] fresh_wire_2058;
	wire [0 : 0] fresh_wire_2059;
	wire [0 : 0] fresh_wire_2060;
	wire [0 : 0] fresh_wire_2061;
	wire [0 : 0] fresh_wire_2062;
	wire [0 : 0] fresh_wire_2063;
	wire [8 : 0] fresh_wire_2064;
	wire [8 : 0] fresh_wire_2065;
	wire [8 : 0] fresh_wire_2066;
	wire [0 : 0] fresh_wire_2067;
	wire [0 : 0] fresh_wire_2068;
	wire [0 : 0] fresh_wire_2069;
	wire [0 : 0] fresh_wire_2070;
	wire [0 : 0] fresh_wire_2071;
	wire [0 : 0] fresh_wire_2072;
	wire [0 : 0] fresh_wire_2073;
	wire [0 : 0] fresh_wire_2074;
	wire [0 : 0] fresh_wire_2075;
	wire [0 : 0] fresh_wire_2076;
	wire [8 : 0] fresh_wire_2077;
	wire [8 : 0] fresh_wire_2078;
	wire [8 : 0] fresh_wire_2079;
	wire [0 : 0] fresh_wire_2080;
	wire [0 : 0] fresh_wire_2081;
	wire [0 : 0] fresh_wire_2082;
	wire [0 : 0] fresh_wire_2083;
	wire [0 : 0] fresh_wire_2084;
	wire [0 : 0] fresh_wire_2085;
	wire [0 : 0] fresh_wire_2086;
	wire [0 : 0] fresh_wire_2087;
	wire [0 : 0] fresh_wire_2088;
	wire [0 : 0] fresh_wire_2089;
	wire [0 : 0] fresh_wire_2090;
	wire [8 : 0] fresh_wire_2091;
	wire [15 : 0] fresh_wire_2092;
	wire [8 : 0] fresh_wire_2093;
	wire [15 : 0] fresh_wire_2094;
	wire [0 : 0] fresh_wire_2095;
	wire [15 : 0] fresh_wire_2096;
	wire [15 : 0] fresh_wire_2097;
	wire [0 : 0] fresh_wire_2098;
	wire [15 : 0] fresh_wire_2099;
	wire [15 : 0] fresh_wire_2100;
	wire [0 : 0] fresh_wire_2101;
	wire [16 : 0] fresh_wire_2102;
	wire [33 : 0] fresh_wire_2103;
	wire [33 : 0] fresh_wire_2104;
	wire [33 : 0] fresh_wire_2105;
	wire [33 : 0] fresh_wire_2106;
	wire [16 : 0] fresh_wire_2107;
	wire [33 : 0] fresh_wire_2108;
	wire [33 : 0] fresh_wire_2109;
	wire [33 : 0] fresh_wire_2110;
	wire [33 : 0] fresh_wire_2111;
	wire [16 : 0] fresh_wire_2112;
	wire [33 : 0] fresh_wire_2113;
	wire [33 : 0] fresh_wire_2114;
	wire [33 : 0] fresh_wire_2115;
	wire [33 : 0] fresh_wire_2116;
	wire [0 : 0] fresh_wire_2117;
	wire [15 : 0] fresh_wire_2118;
	wire [16 : 0] fresh_wire_2119;
	wire [15 : 0] fresh_wire_2120;
	wire [16 : 0] fresh_wire_2121;
	wire [16 : 0] fresh_wire_2122;
	wire [16 : 0] fresh_wire_2123;
	wire [16 : 0] fresh_wire_2124;
	wire [16 : 0] fresh_wire_2125;
	wire [16 : 0] fresh_wire_2126;
	wire [16 : 0] fresh_wire_2127;
	wire [15 : 0] fresh_wire_2128;
	wire [16 : 0] fresh_wire_2129;
	wire [15 : 0] fresh_wire_2130;
	wire [16 : 0] fresh_wire_2131;
	wire [16 : 0] fresh_wire_2132;
	wire [16 : 0] fresh_wire_2133;
	wire [16 : 0] fresh_wire_2134;
	wire [16 : 0] fresh_wire_2135;
	wire [16 : 0] fresh_wire_2136;
	wire [16 : 0] fresh_wire_2137;
	wire [16 : 0] fresh_wire_2138;
	wire [33 : 0] fresh_wire_2139;
	wire [33 : 0] fresh_wire_2140;
	wire [33 : 0] fresh_wire_2141;
	wire [33 : 0] fresh_wire_2142;
	wire [15 : 0] fresh_wire_2143;
	wire [15 : 0] fresh_wire_2144;
	wire [0 : 0] fresh_wire_2145;
	wire [0 : 0] fresh_wire_2146;
	wire [16 : 0] fresh_wire_2147;
	wire [33 : 0] fresh_wire_2148;
	wire [33 : 0] fresh_wire_2149;
	wire [33 : 0] fresh_wire_2150;
	wire [33 : 0] fresh_wire_2151;
	wire [15 : 0] fresh_wire_2152;
	wire [16 : 0] fresh_wire_2153;
	wire [15 : 0] fresh_wire_2154;
	wire [16 : 0] fresh_wire_2155;
	wire [16 : 0] fresh_wire_2156;
	wire [16 : 0] fresh_wire_2157;
	wire [16 : 0] fresh_wire_2158;
	wire [16 : 0] fresh_wire_2159;
	wire [16 : 0] fresh_wire_2160;
	wire [16 : 0] fresh_wire_2161;
	wire [15 : 0] fresh_wire_2162;
	wire [16 : 0] fresh_wire_2163;
	wire [15 : 0] fresh_wire_2164;
	wire [16 : 0] fresh_wire_2165;
	wire [16 : 0] fresh_wire_2166;
	wire [16 : 0] fresh_wire_2167;
	wire [16 : 0] fresh_wire_2168;
	wire [16 : 0] fresh_wire_2169;
	wire [16 : 0] fresh_wire_2170;
	wire [16 : 0] fresh_wire_2171;
	wire [16 : 0] fresh_wire_2172;
	wire [33 : 0] fresh_wire_2173;
	wire [33 : 0] fresh_wire_2174;
	wire [33 : 0] fresh_wire_2175;
	wire [33 : 0] fresh_wire_2176;
	wire [0 : 0] fresh_wire_2177;
	wire [15 : 0] fresh_wire_2178;
	wire [16 : 0] fresh_wire_2179;
	wire [16 : 0] fresh_wire_2180;
	wire [16 : 0] fresh_wire_2181;
	wire [16 : 0] fresh_wire_2182;
	wire [16 : 0] fresh_wire_2183;
	wire [16 : 0] fresh_wire_2184;
	wire [16 : 0] fresh_wire_2185;
	wire [15 : 0] fresh_wire_2186;
	wire [16 : 0] fresh_wire_2187;
	wire [15 : 0] fresh_wire_2188;
	wire [16 : 0] fresh_wire_2189;
	wire [16 : 0] fresh_wire_2190;
	wire [16 : 0] fresh_wire_2191;
	wire [16 : 0] fresh_wire_2192;
	wire [16 : 0] fresh_wire_2193;
	wire [16 : 0] fresh_wire_2194;
	wire [16 : 0] fresh_wire_2195;
	wire [15 : 0] fresh_wire_2196;
	wire [16 : 0] fresh_wire_2197;
	wire [15 : 0] fresh_wire_2198;
	wire [16 : 0] fresh_wire_2199;
	wire [16 : 0] fresh_wire_2200;
	wire [16 : 0] fresh_wire_2201;
	wire [16 : 0] fresh_wire_2202;
	wire [16 : 0] fresh_wire_2203;
	wire [16 : 0] fresh_wire_2204;
	wire [16 : 0] fresh_wire_2205;
	wire [15 : 0] fresh_wire_2206;
	wire [16 : 0] fresh_wire_2207;
	wire [15 : 0] fresh_wire_2208;
	wire [16 : 0] fresh_wire_2209;
	wire [16 : 0] fresh_wire_2210;
	wire [16 : 0] fresh_wire_2211;
	wire [16 : 0] fresh_wire_2212;
	wire [16 : 0] fresh_wire_2213;
	wire [16 : 0] fresh_wire_2214;
	wire [16 : 0] fresh_wire_2215;
	wire [16 : 0] fresh_wire_2216;
	wire [33 : 0] fresh_wire_2217;
	wire [33 : 0] fresh_wire_2218;
	wire [33 : 0] fresh_wire_2219;
	wire [33 : 0] fresh_wire_2220;
	wire [15 : 0] fresh_wire_2221;
	wire [15 : 0] fresh_wire_2222;
	wire [0 : 0] fresh_wire_2223;
	wire [0 : 0] fresh_wire_2224;
	wire [16 : 0] fresh_wire_2225;
	wire [33 : 0] fresh_wire_2226;
	wire [33 : 0] fresh_wire_2227;
	wire [33 : 0] fresh_wire_2228;
	wire [33 : 0] fresh_wire_2229;
	wire [15 : 0] fresh_wire_2230;
	wire [15 : 0] fresh_wire_2231;
	wire [0 : 0] fresh_wire_2232;
	wire [0 : 0] fresh_wire_2233;
	wire [16 : 0] fresh_wire_2234;
	wire [33 : 0] fresh_wire_2235;
	wire [33 : 0] fresh_wire_2236;
	wire [33 : 0] fresh_wire_2237;
	wire [33 : 0] fresh_wire_2238;
	wire [15 : 0] fresh_wire_2239;
	wire [16 : 0] fresh_wire_2240;
	wire [15 : 0] fresh_wire_2241;
	wire [16 : 0] fresh_wire_2242;
	wire [16 : 0] fresh_wire_2243;
	wire [16 : 0] fresh_wire_2244;
	wire [16 : 0] fresh_wire_2245;
	wire [16 : 0] fresh_wire_2246;
	wire [16 : 0] fresh_wire_2247;
	wire [16 : 0] fresh_wire_2248;
	wire [0 : 0] fresh_wire_2249;
	wire [0 : 0] fresh_wire_2250;
	wire [15 : 0] fresh_wire_2251;
	wire [15 : 0] fresh_wire_2252;
	wire [15 : 0] fresh_wire_2253;
	wire [15 : 0] fresh_wire_2254;
	wire [15 : 0] fresh_wire_2255;
	wire [15 : 0] fresh_wire_2256;
	wire [15 : 0] fresh_wire_2257;
	wire [15 : 0] fresh_wire_2258;
	wire [15 : 0] fresh_wire_2259;
	wire [15 : 0] fresh_wire_2260;
	wire [15 : 0] fresh_wire_2261;
	wire [15 : 0] fresh_wire_2262;
	wire [15 : 0] fresh_wire_2263;
	wire [15 : 0] fresh_wire_2264;
	wire [15 : 0] fresh_wire_2265;
	wire [15 : 0] fresh_wire_2266;
	wire [15 : 0] fresh_wire_2267;
	wire [15 : 0] fresh_wire_2268;
	wire [0 : 0] fresh_wire_2269;
	wire [33 : 0] fresh_wire_2270;
	wire [0 : 0] fresh_wire_2271;
	wire [33 : 0] fresh_wire_2272;
	wire [0 : 0] fresh_wire_2273;
	wire [33 : 0] fresh_wire_2274;
	wire [0 : 0] fresh_wire_2275;
	wire [0 : 0] fresh_wire_2276;
	wire [0 : 0] fresh_wire_2277;
	wire [0 : 0] fresh_wire_2278;
	wire [16 : 0] fresh_wire_2279;
	wire [16 : 0] fresh_wire_2280;
	wire [0 : 0] fresh_wire_2281;
	wire [33 : 0] fresh_wire_2282;
	wire [0 : 0] fresh_wire_2283;
	wire [0 : 0] fresh_wire_2284;
	wire [33 : 0] fresh_wire_2285;
	wire [16 : 0] fresh_wire_2286;
	wire [16 : 0] fresh_wire_2287;
	wire [0 : 0] fresh_wire_2288;
	wire [33 : 0] fresh_wire_2289;
	wire [0 : 0] fresh_wire_2290;
	wire [0 : 0] fresh_wire_2291;
	wire [0 : 0] fresh_wire_2292;
	wire [0 : 0] fresh_wire_2293;
	wire [16 : 0] fresh_wire_2294;
	wire [16 : 0] fresh_wire_2295;
	wire [16 : 0] fresh_wire_2296;
	wire [16 : 0] fresh_wire_2297;
	wire [16 : 0] fresh_wire_2298;
	wire [0 : 0] fresh_wire_2299;
	wire [33 : 0] fresh_wire_2300;
	wire [0 : 0] fresh_wire_2301;
	wire [0 : 0] fresh_wire_2302;
	wire [33 : 0] fresh_wire_2303;
	wire [0 : 0] fresh_wire_2304;
	wire [0 : 0] fresh_wire_2305;
	wire [33 : 0] fresh_wire_2306;
	wire [16 : 0] fresh_wire_2307;
	wire [0 : 0] fresh_wire_2308;
	wire [0 : 0] fresh_wire_2309;
	wire [0 : 0] fresh_wire_2310;
	wire [0 : 0] fresh_wire_2311;
	wire [0 : 0] fresh_wire_2312;
	wire [0 : 0] fresh_wire_2313;
	wire [0 : 0] fresh_wire_2314;
	wire [0 : 0] fresh_wire_2315;
	wire [0 : 0] fresh_wire_2316;
	wire [0 : 0] fresh_wire_2317;
	wire [0 : 0] fresh_wire_2318;
	wire [0 : 0] fresh_wire_2319;
	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) aux_div_pad_port_cell(.PORT_ID_IN(fresh_wire_0),
.PORT_ID_OUT(aux_div_pad));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) cell_149_3_const_replacement(.PORT_ID_OUT(fresh_wire_2250));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) cell_261940_3_const_replacement(.PORT_ID_OUT(fresh_wire_2269));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(34'h000000013),
.PARAM_WIDTH(32'h00000022)) cell_261945_3_const_replacement(.PORT_ID_OUT(fresh_wire_2270));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(16'h0001),
.PARAM_WIDTH(32'h00000010)) cell_26382_3_const_replacement(.PORT_ID_OUT(fresh_wire_2251));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(16'h0002),
.PARAM_WIDTH(32'h00000010)) cell_26400_3_const_replacement(.PORT_ID_OUT(fresh_wire_2252));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(16'h0002),
.PARAM_WIDTH(32'h00000010)) cell_26409_3_const_replacement(.PORT_ID_OUT(fresh_wire_2253));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(16'h0001),
.PARAM_WIDTH(32'h00000010)) cell_26415_3_const_replacement(.PORT_ID_OUT(fresh_wire_2254));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(16'h0040),
.PARAM_WIDTH(32'h00000010)) cell_26436_3_const_replacement(.PORT_ID_OUT(fresh_wire_2255));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) cell_264628_3_const_replacement(.PORT_ID_OUT(fresh_wire_2271));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(34'h000000010),
.PARAM_WIDTH(32'h00000022)) cell_264633_3_const_replacement(.PORT_ID_OUT(fresh_wire_2272));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(16'h0040),
.PARAM_WIDTH(32'h00000010)) cell_26550_3_const_replacement(.PORT_ID_OUT(fresh_wire_2256));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_26608_3_const_replacement(.PORT_ID_OUT(fresh_wire_2308));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_26618_3_const_replacement(.PORT_ID_OUT(fresh_wire_2309));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_26641_3_const_replacement(.PORT_ID_OUT(fresh_wire_2310));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_26648_3_const_replacement(.PORT_ID_OUT(fresh_wire_2311));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_26668_3_const_replacement(.PORT_ID_OUT(fresh_wire_2312));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) cell_26671_3_const_replacement(.PORT_ID_OUT(fresh_wire_2313));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) cell_267321_3_const_replacement(.PORT_ID_OUT(fresh_wire_2273));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(34'h000000012),
.PARAM_WIDTH(32'h00000022)) cell_267326_3_const_replacement(.PORT_ID_OUT(fresh_wire_2274));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(16'h0040),
.PARAM_WIDTH(32'h00000010)) cell_26849_3_const_replacement(.PORT_ID_OUT(fresh_wire_2257));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(16'h001f),
.PARAM_WIDTH(32'h00000010)) cell_26860_3_const_replacement(.PORT_ID_OUT(fresh_wire_2258));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(16'h003b),
.PARAM_WIDTH(32'h00000010)) cell_26866_3_const_replacement(.PORT_ID_OUT(fresh_wire_2259));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_27034_3_const_replacement(.PORT_ID_OUT(fresh_wire_2275));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_27039_3_const_replacement(.PORT_ID_OUT(fresh_wire_2276));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_27064_3_const_replacement(.PORT_ID_OUT(fresh_wire_2277));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_27069_3_const_replacement(.PORT_ID_OUT(fresh_wire_2278));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(17'h00000),
.PARAM_WIDTH(32'h00000011)) cell_293878_3_const_replacement(.PORT_ID_OUT(fresh_wire_2279));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(17'h00000),
.PARAM_WIDTH(32'h00000011)) cell_296571_3_const_replacement(.PORT_ID_OUT(fresh_wire_2280));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) cell_299632_3_const_replacement(.PORT_ID_OUT(fresh_wire_2281));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(34'h000000000),
.PARAM_WIDTH(32'h00000022)) cell_299637_3_const_replacement(.PORT_ID_OUT(fresh_wire_2282));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_299833_3_const_replacement(.PORT_ID_OUT(fresh_wire_2283));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) cell_302320_3_const_replacement(.PORT_ID_OUT(fresh_wire_2284));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(34'h00000000c),
.PARAM_WIDTH(32'h00000022)) cell_302325_3_const_replacement(.PORT_ID_OUT(fresh_wire_2285));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(17'h00000),
.PARAM_WIDTH(32'h00000011)) cell_326139_3_const_replacement(.PORT_ID_OUT(fresh_wire_2286));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(17'h00000),
.PARAM_WIDTH(32'h00000011)) cell_328832_3_const_replacement(.PORT_ID_OUT(fresh_wire_2287));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) cell_331893_3_const_replacement(.PORT_ID_OUT(fresh_wire_2288));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(34'h000000011),
.PARAM_WIDTH(32'h00000022)) cell_331898_3_const_replacement(.PORT_ID_OUT(fresh_wire_2289));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(17'h00000),
.PARAM_WIDTH(32'h00000011)) cell_336893_3_const_replacement(.PORT_ID_OUT(fresh_wire_2295));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(17'h00000),
.PARAM_WIDTH(32'h00000011)) cell_336896_3_const_replacement(.PORT_ID_OUT(fresh_wire_2294));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(17'h00000),
.PARAM_WIDTH(32'h00000011)) cell_358400_3_const_replacement(.PORT_ID_OUT(fresh_wire_2296));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(17'h00000),
.PARAM_WIDTH(32'h00000011)) cell_361093_3_const_replacement(.PORT_ID_OUT(fresh_wire_2297));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(17'h00000),
.PARAM_WIDTH(32'h00000011)) cell_363781_3_const_replacement(.PORT_ID_OUT(fresh_wire_2298));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) cell_366842_3_const_replacement(.PORT_ID_OUT(fresh_wire_2299));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(34'h00000000e),
.PARAM_WIDTH(32'h00000022)) cell_366847_3_const_replacement(.PORT_ID_OUT(fresh_wire_2300));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_367043_3_const_replacement(.PORT_ID_OUT(fresh_wire_2301));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) cell_369530_3_const_replacement(.PORT_ID_OUT(fresh_wire_2302));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(34'h00000000b),
.PARAM_WIDTH(32'h00000022)) cell_369535_3_const_replacement(.PORT_ID_OUT(fresh_wire_2303));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_391240_3_const_replacement(.PORT_ID_OUT(fresh_wire_2304));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) cell_393727_3_const_replacement(.PORT_ID_OUT(fresh_wire_2305));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(34'h00000000d),
.PARAM_WIDTH(32'h00000022)) cell_393732_3_const_replacement(.PORT_ID_OUT(fresh_wire_2306));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(17'h00000),
.PARAM_WIDTH(32'h00000011)) cell_398730_3_const_replacement(.PORT_ID_OUT(fresh_wire_2307));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(16'h0001),
.PARAM_WIDTH(32'h00000010)) cell_52015_3_const_replacement(.PORT_ID_OUT(fresh_wire_2260));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(16'h0002),
.PARAM_WIDTH(32'h00000010)) cell_52033_3_const_replacement(.PORT_ID_OUT(fresh_wire_2261));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(16'h0002),
.PARAM_WIDTH(32'h00000010)) cell_52042_3_const_replacement(.PORT_ID_OUT(fresh_wire_2262));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(16'h0001),
.PARAM_WIDTH(32'h00000010)) cell_52048_3_const_replacement(.PORT_ID_OUT(fresh_wire_2263));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(16'h0040),
.PARAM_WIDTH(32'h00000010)) cell_52069_3_const_replacement(.PORT_ID_OUT(fresh_wire_2264));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(16'h0040),
.PARAM_WIDTH(32'h00000010)) cell_52183_3_const_replacement(.PORT_ID_OUT(fresh_wire_2265));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_52241_3_const_replacement(.PORT_ID_OUT(fresh_wire_2314));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_52251_3_const_replacement(.PORT_ID_OUT(fresh_wire_2315));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_52274_3_const_replacement(.PORT_ID_OUT(fresh_wire_2316));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_52281_3_const_replacement(.PORT_ID_OUT(fresh_wire_2317));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_52301_3_const_replacement(.PORT_ID_OUT(fresh_wire_2318));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) cell_52304_3_const_replacement(.PORT_ID_OUT(fresh_wire_2319));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(16'h0040),
.PARAM_WIDTH(32'h00000010)) cell_52482_3_const_replacement(.PORT_ID_OUT(fresh_wire_2266));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(16'h001f),
.PARAM_WIDTH(32'h00000010)) cell_52493_3_const_replacement(.PORT_ID_OUT(fresh_wire_2267));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(16'h003b),
.PARAM_WIDTH(32'h00000010)) cell_52499_3_const_replacement(.PORT_ID_OUT(fresh_wire_2268));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_52667_3_const_replacement(.PORT_ID_OUT(fresh_wire_2290));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_52672_3_const_replacement(.PORT_ID_OUT(fresh_wire_2291));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_52697_3_const_replacement(.PORT_ID_OUT(fresh_wire_2292));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) cell_52702_3_const_replacement(.PORT_ID_OUT(fresh_wire_2293));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) clk_ext_in_port_cell(.PORT_ID_IN(clk_ext_in),
.PORT_ID_OUT(fresh_wire_1));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) clk_in_port_cell(.PORT_ID_IN(clk_in),
.PORT_ID_OUT(fresh_wire_2));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000020),
.PARAM_PORT_TYPE(2'h0)) config_addr_in_port_cell(.PORT_ID_IN(config_addr_in),
.PORT_ID_OUT(fresh_wire_3));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000020),
.PARAM_PORT_TYPE(2'h0)) config_data_in_port_cell(.PORT_ID_IN(config_data_in),
.PORT_ID_OUT(fresh_wire_4));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) ext_cki_jm_port_cell(.PORT_ID_IN(ext_cki_jm),
.PORT_ID_OUT(fresh_wire_6));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) ext_cki_port_cell(.PORT_ID_IN(ext_cki),
.PORT_ID_OUT(fresh_wire_5));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) ext_ckib_jm_port_cell(.PORT_ID_IN(ext_ckib_jm),
.PORT_ID_OUT(fresh_wire_8));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) ext_ckib_port_cell(.PORT_ID_IN(ext_ckib),
.PORT_ID_OUT(fresh_wire_7));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) ext_frefn_jm_port_cell(.PORT_ID_IN(ext_frefn_jm),
.PORT_ID_OUT(fresh_wire_10));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) ext_frefn_port_cell(.PORT_ID_IN(ext_frefn),
.PORT_ID_OUT(fresh_wire_9));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) ext_frefp_jm_port_cell(.PORT_ID_IN(ext_frefp_jm),
.PORT_ID_OUT(fresh_wire_12));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) ext_frefp_port_cell(.PORT_ID_IN(ext_frefp),
.PORT_ID_OUT(fresh_wire_11));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) ffeed_pad_port_cell(.PORT_ID_IN(fresh_wire_13),
.PORT_ID_OUT(ffeed_pad));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) fout_div_pad_port_cell(.PORT_ID_IN(fresh_wire_14),
.PORT_ID_OUT(fout_div_pad));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) fref_off_pad_port_cell(.PORT_ID_IN(fresh_wire_15),
.PORT_ID_OUT(fref_off_pad));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) frefn_out_jm_port_cell(.PORT_ID_IN(fresh_wire_16),
.PORT_ID_OUT(frefn_out_jm));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) frefp_out_jm_port_cell(.PORT_ID_IN(fresh_wire_17),
.PORT_ID_OUT(frefp_out_jm));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h0000000d),
.PARAM_PORT_TYPE(2'h1)) lf_out_port_cell(.PORT_ID_IN(fresh_wire_18),
.PORT_ID_OUT(lf_out));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(13'h0000),
.PARAM_WIDTH(32'h0000000d)) mdll_top$self_lf_out(.PORT_ID_OUT(fresh_wire_154));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000004),
.PARAM_PORT_TYPE(2'h1)) mdllout_pad_port_cell(.PORT_ID_IN(fresh_wire_19),
.PORT_ID_OUT(mdllout_pad));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$__DOLLAR__and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__memory_core_unq1__DOT__v__COLON__309__DOLLAR__631$op0(.PORT_ID_IN0(fresh_wire_155),
.PORT_ID_IN1(fresh_wire_156),
.PORT_ID_OUT(fresh_wire_157));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$__DOLLAR__and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__memory_core_unq1__DOT__v__COLON__310__DOLLAR__633$op0(.PORT_ID_IN0(fresh_wire_158),
.PORT_ID_IN1(fresh_wire_159),
.PORT_ID_OUT(fresh_wire_160));

	CELL_TYPE_OR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$__DOLLAR__or__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__memory_core_unq1__DOT__v__COLON__309__DOLLAR__630$op0(.PORT_ID_IN0(fresh_wire_161),
.PORT_ID_IN1(fresh_wire_162),
.PORT_ID_OUT(fresh_wire_163));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__471$op0(.PORT_ID_IN0(fresh_wire_164),
.PORT_ID_IN1(fresh_wire_165),
.PORT_ID_OUT(fresh_wire_166));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000002),
.PARAM_OUT_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__206__DOLLAR__488$extendB(.PORT_ID_IN(fresh_wire_167),
.PORT_ID_OUT(fresh_wire_168));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__206__DOLLAR__488$op0(.PORT_ID_IN0(fresh_wire_169),
.PORT_ID_IN1(fresh_wire_170),
.PORT_ID_OUT(fresh_wire_171));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__233__DOLLAR__500$extendA(.PORT_ID_IN(fresh_wire_172),
.PORT_ID_OUT(fresh_wire_173));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__233__DOLLAR__500$op0(.PORT_ID_IN0(fresh_wire_174),
.PORT_ID_IN1(fresh_wire_175),
.PORT_ID_OUT(fresh_wire_176));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__235__DOLLAR__501$extendA(.PORT_ID_IN(fresh_wire_177),
.PORT_ID_OUT(fresh_wire_178));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__235__DOLLAR__501$op0(.PORT_ID_IN0(fresh_wire_179),
.PORT_ID_IN1(fresh_wire_180),
.PORT_ID_OUT(fresh_wire_181));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__242__DOLLAR__504$extendA(.PORT_ID_IN(fresh_wire_182),
.PORT_ID_OUT(fresh_wire_183));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__242__DOLLAR__504$op0(.PORT_ID_IN0(fresh_wire_184),
.PORT_ID_IN1(fresh_wire_185),
.PORT_ID_OUT(fresh_wire_186));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__271__DOLLAR__521$op0(.PORT_ID_IN0(fresh_wire_187),
.PORT_ID_IN1(fresh_wire_188),
.PORT_ID_OUT(fresh_wire_189));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__273__DOLLAR__525$op0(.PORT_ID_IN0(fresh_wire_190),
.PORT_ID_IN1(fresh_wire_191),
.PORT_ID_OUT(fresh_wire_192));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__276__DOLLAR__534$op0(.PORT_ID_IN0(fresh_wire_193),
.PORT_ID_IN1(fresh_wire_194),
.PORT_ID_OUT(fresh_wire_195));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__555$op0(.PORT_ID_IN0(fresh_wire_196),
.PORT_ID_IN1(fresh_wire_197),
.PORT_ID_OUT(fresh_wire_198));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__207__DOLLAR__491$op0(.PORT_ID_IN0(fresh_wire_199),
.PORT_ID_IN1(fresh_wire_200),
.PORT_ID_OUT(fresh_wire_201));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__466$op0(.PORT_ID_IN0(fresh_wire_202),
.PORT_ID_IN1(fresh_wire_203),
.PORT_ID_OUT(fresh_wire_204));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__467$op0(.PORT_ID_IN0(fresh_wire_205),
.PORT_ID_IN1(fresh_wire_206),
.PORT_ID_OUT(fresh_wire_207));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__469$op0(.PORT_ID_IN0(fresh_wire_208),
.PORT_ID_IN1(fresh_wire_209),
.PORT_ID_OUT(fresh_wire_210));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__472$op0(.PORT_ID_IN0(fresh_wire_211),
.PORT_ID_IN1(fresh_wire_212),
.PORT_ID_OUT(fresh_wire_213));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__176__DOLLAR__474$op0(.PORT_ID_IN0(fresh_wire_214),
.PORT_ID_IN1(fresh_wire_215),
.PORT_ID_OUT(fresh_wire_216));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__192__DOLLAR__482$op0(.PORT_ID_IN0(fresh_wire_217),
.PORT_ID_IN1(fresh_wire_218),
.PORT_ID_OUT(fresh_wire_219));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__193__DOLLAR__483$op0(.PORT_ID_IN0(fresh_wire_220),
.PORT_ID_IN1(fresh_wire_221),
.PORT_ID_OUT(fresh_wire_222));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__196__DOLLAR__484$op0(.PORT_ID_IN0(fresh_wire_223),
.PORT_ID_IN1(fresh_wire_224),
.PORT_ID_OUT(fresh_wire_225));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__207__DOLLAR__490$op0(.PORT_ID_IN0(fresh_wire_226),
.PORT_ID_IN1(fresh_wire_227),
.PORT_ID_OUT(fresh_wire_228));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__228__DOLLAR__497$op0(.PORT_ID_IN0(fresh_wire_229),
.PORT_ID_IN1(fresh_wire_230),
.PORT_ID_OUT(fresh_wire_231));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__229__DOLLAR__498$op0(.PORT_ID_IN0(fresh_wire_232),
.PORT_ID_IN1(fresh_wire_233),
.PORT_ID_OUT(fresh_wire_234));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__268__DOLLAR__513$op0(.PORT_ID_IN0(fresh_wire_235),
.PORT_ID_IN1(fresh_wire_236),
.PORT_ID_OUT(fresh_wire_237));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__268__DOLLAR__516$op0(.PORT_ID_IN0(fresh_wire_238),
.PORT_ID_IN1(fresh_wire_239),
.PORT_ID_OUT(fresh_wire_240));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__273__DOLLAR__524$op0(.PORT_ID_IN0(fresh_wire_241),
.PORT_ID_IN1(fresh_wire_242),
.PORT_ID_OUT(fresh_wire_243));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__285__DOLLAR__541$op0(.PORT_ID_IN0(fresh_wire_244),
.PORT_ID_IN1(fresh_wire_245),
.PORT_ID_OUT(fresh_wire_246));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__309__DOLLAR__549$op0(.PORT_ID_IN0(fresh_wire_247),
.PORT_ID_IN1(fresh_wire_248),
.PORT_ID_OUT(fresh_wire_249));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__556$op0(.PORT_ID_IN0(fresh_wire_250),
.PORT_ID_IN1(fresh_wire_251),
.PORT_ID_OUT(fresh_wire_252));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__316__DOLLAR__558$op0(.PORT_ID_IN0(fresh_wire_253),
.PORT_ID_IN1(fresh_wire_254),
.PORT_ID_OUT(fresh_wire_255));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__355__DOLLAR__568$op0(.PORT_ID_IN0(fresh_wire_256),
.PORT_ID_IN1(fresh_wire_257),
.PORT_ID_OUT(fresh_wire_258));

	CELL_TYPE_UGE #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__ge__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__230__DOLLAR__499$op0(.PORT_ID_IN0(fresh_wire_259),
.PORT_ID_IN1(fresh_wire_260),
.PORT_ID_OUT(fresh_wire_261));

	CELL_TYPE_UGE #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__ge__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__239__DOLLAR__503$op0(.PORT_ID_IN0(fresh_wire_262),
.PORT_ID_IN1(fresh_wire_263),
.PORT_ID_OUT(fresh_wire_264));

	CELL_TYPE_UGE #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__ge__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__276__DOLLAR__535$op0(.PORT_ID_IN0(fresh_wire_265),
.PORT_ID_IN1(fresh_wire_266),
.PORT_ID_OUT(fresh_wire_267));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__468$aRed(.PORT_ID_IN(fresh_wire_268),
.PORT_ID_OUT(fresh_wire_269));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__468$andOps(.PORT_ID_IN0(fresh_wire_270),
.PORT_ID_IN1(fresh_wire_271),
.PORT_ID_OUT(fresh_wire_272));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__468$bRed(.PORT_ID_IN(fresh_wire_273),
.PORT_ID_OUT(fresh_wire_274));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__470$aRed(.PORT_ID_IN(fresh_wire_275),
.PORT_ID_OUT(fresh_wire_276));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__470$andOps(.PORT_ID_IN0(fresh_wire_277),
.PORT_ID_IN1(fresh_wire_278),
.PORT_ID_OUT(fresh_wire_279));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__470$bRed(.PORT_ID_IN(fresh_wire_280),
.PORT_ID_OUT(fresh_wire_281));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__473$aRed(.PORT_ID_IN(fresh_wire_282),
.PORT_ID_OUT(fresh_wire_283));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__473$andOps(.PORT_ID_IN0(fresh_wire_284),
.PORT_ID_IN1(fresh_wire_285),
.PORT_ID_OUT(fresh_wire_286));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__473$bRed(.PORT_ID_IN(fresh_wire_287),
.PORT_ID_OUT(fresh_wire_288));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__268__DOLLAR__515$aRed(.PORT_ID_IN(fresh_wire_289),
.PORT_ID_OUT(fresh_wire_290));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__268__DOLLAR__515$andOps(.PORT_ID_IN0(fresh_wire_291),
.PORT_ID_IN1(fresh_wire_292),
.PORT_ID_OUT(fresh_wire_293));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__268__DOLLAR__517$aRed(.PORT_ID_IN(fresh_wire_294),
.PORT_ID_OUT(fresh_wire_295));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__268__DOLLAR__517$andOps(.PORT_ID_IN0(fresh_wire_296),
.PORT_ID_IN1(fresh_wire_297),
.PORT_ID_OUT(fresh_wire_298));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__268__DOLLAR__517$bRed(.PORT_ID_IN(fresh_wire_299),
.PORT_ID_OUT(fresh_wire_300));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__271__DOLLAR__520$aRed(.PORT_ID_IN(fresh_wire_301),
.PORT_ID_OUT(fresh_wire_302));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__271__DOLLAR__520$andOps(.PORT_ID_IN0(fresh_wire_303),
.PORT_ID_IN1(fresh_wire_304),
.PORT_ID_OUT(fresh_wire_305));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__271__DOLLAR__523$aRed(.PORT_ID_IN(fresh_wire_306),
.PORT_ID_OUT(fresh_wire_307));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__271__DOLLAR__523$andOps(.PORT_ID_IN0(fresh_wire_308),
.PORT_ID_IN1(fresh_wire_309),
.PORT_ID_OUT(fresh_wire_310));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__271__DOLLAR__523$bRed(.PORT_ID_IN(fresh_wire_311),
.PORT_ID_OUT(fresh_wire_312));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__276__DOLLAR__536$aRed(.PORT_ID_IN(fresh_wire_313),
.PORT_ID_OUT(fresh_wire_314));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__276__DOLLAR__536$andOps(.PORT_ID_IN0(fresh_wire_315),
.PORT_ID_IN1(fresh_wire_316),
.PORT_ID_OUT(fresh_wire_317));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__276__DOLLAR__536$bRed(.PORT_ID_IN(fresh_wire_318),
.PORT_ID_OUT(fresh_wire_319));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__277__DOLLAR__539$andOps(.PORT_ID_IN0(fresh_wire_320),
.PORT_ID_IN1(fresh_wire_321),
.PORT_ID_OUT(fresh_wire_322));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__277__DOLLAR__539$bRed(.PORT_ID_IN(fresh_wire_323),
.PORT_ID_OUT(fresh_wire_324));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__285__DOLLAR__543$aRed(.PORT_ID_IN(fresh_wire_325),
.PORT_ID_OUT(fresh_wire_326));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__285__DOLLAR__543$andOps(.PORT_ID_IN0(fresh_wire_327),
.PORT_ID_IN1(fresh_wire_328),
.PORT_ID_OUT(fresh_wire_329));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__552$aRed(.PORT_ID_IN(fresh_wire_330),
.PORT_ID_OUT(fresh_wire_331));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__552$andOps(.PORT_ID_IN0(fresh_wire_332),
.PORT_ID_IN1(fresh_wire_333),
.PORT_ID_OUT(fresh_wire_334));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__552$bRed(.PORT_ID_IN(fresh_wire_335),
.PORT_ID_OUT(fresh_wire_336));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__554$aRed(.PORT_ID_IN(fresh_wire_337),
.PORT_ID_OUT(fresh_wire_338));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__554$andOps(.PORT_ID_IN0(fresh_wire_339),
.PORT_ID_IN1(fresh_wire_340),
.PORT_ID_OUT(fresh_wire_341));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__554$bRed(.PORT_ID_IN(fresh_wire_342),
.PORT_ID_OUT(fresh_wire_343));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__557$aRed(.PORT_ID_IN(fresh_wire_344),
.PORT_ID_OUT(fresh_wire_345));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__557$andOps(.PORT_ID_IN0(fresh_wire_346),
.PORT_ID_IN1(fresh_wire_347),
.PORT_ID_OUT(fresh_wire_348));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__557$bRed(.PORT_ID_IN(fresh_wire_349),
.PORT_ID_OUT(fresh_wire_350));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__316__DOLLAR__560$aRed(.PORT_ID_IN(fresh_wire_351),
.PORT_ID_OUT(fresh_wire_352));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__316__DOLLAR__560$andOps(.PORT_ID_IN0(fresh_wire_353),
.PORT_ID_IN1(fresh_wire_354),
.PORT_ID_OUT(fresh_wire_355));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_or__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__344__DOLLAR__565$bRed(.PORT_ID_IN(fresh_wire_356),
.PORT_ID_OUT(fresh_wire_357));

	CELL_TYPE_OR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__logic_or__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__344__DOLLAR__565$orOps(.PORT_ID_IN0(fresh_wire_358),
.PORT_ID_IN1(fresh_wire_359),
.PORT_ID_OUT(fresh_wire_360));

	CELL_TYPE_ULT #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__lt__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__250__DOLLAR__507$op0(.PORT_ID_IN0(fresh_wire_361),
.PORT_ID_IN1(fresh_wire_362),
.PORT_ID_OUT(fresh_wire_363));

	CELL_TYPE_ULT #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__lt__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__271__DOLLAR__522$op0(.PORT_ID_IN0(fresh_wire_364),
.PORT_ID_IN1(fresh_wire_365),
.PORT_ID_OUT(fresh_wire_366));

	CELL_TYPE_NOT #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__not__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__171__DOLLAR__465$op0(.PORT_ID_IN(fresh_wire_367),
.PORT_ID_OUT(fresh_wire_368));

	CELL_TYPE_REG #(.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3712$reg0(.PORT_ID_CLK(fresh_wire_371),
.PORT_ID_IN(fresh_wire_369),
.PORT_ID_OUT(fresh_wire_370));

	CELL_TYPE_REG #(.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(2'hx),
.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3713$reg0(.PORT_ID_CLK(fresh_wire_374),
.PORT_ID_IN(fresh_wire_372),
.PORT_ID_OUT(fresh_wire_373));

	CELL_TYPE_REG #(.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(2'hx),
.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3714$reg0(.PORT_ID_CLK(fresh_wire_377),
.PORT_ID_IN(fresh_wire_375),
.PORT_ID_OUT(fresh_wire_376));

	CELL_TYPE_REG #(.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(16'hxxxx),
.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3716$reg0(.PORT_ID_CLK(fresh_wire_380),
.PORT_ID_IN(fresh_wire_378),
.PORT_ID_OUT(fresh_wire_379));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3718$reg0(.PORT_ID_ARST(fresh_wire_384),
.PORT_ID_CLK(fresh_wire_383),
.PORT_ID_IN(fresh_wire_381),
.PORT_ID_OUT(fresh_wire_382));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3719$reg0(.PORT_ID_ARST(fresh_wire_388),
.PORT_ID_CLK(fresh_wire_387),
.PORT_ID_IN(fresh_wire_385),
.PORT_ID_OUT(fresh_wire_386));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3720$reg0(.PORT_ID_ARST(fresh_wire_392),
.PORT_ID_CLK(fresh_wire_391),
.PORT_ID_IN(fresh_wire_389),
.PORT_ID_OUT(fresh_wire_390));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3721$reg0(.PORT_ID_ARST(fresh_wire_396),
.PORT_ID_CLK(fresh_wire_395),
.PORT_ID_IN(fresh_wire_393),
.PORT_ID_OUT(fresh_wire_394));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3722$reg0(.PORT_ID_ARST(fresh_wire_400),
.PORT_ID_CLK(fresh_wire_399),
.PORT_ID_IN(fresh_wire_397),
.PORT_ID_OUT(fresh_wire_398));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(2'h0),
.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3723$reg0(.PORT_ID_ARST(fresh_wire_404),
.PORT_ID_CLK(fresh_wire_403),
.PORT_ID_IN(fresh_wire_401),
.PORT_ID_OUT(fresh_wire_402));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(16'h0000),
.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3724$reg0(.PORT_ID_ARST(fresh_wire_408),
.PORT_ID_CLK(fresh_wire_407),
.PORT_ID_IN(fresh_wire_405),
.PORT_ID_OUT(fresh_wire_406));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(16'h0000),
.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3725$reg0(.PORT_ID_ARST(fresh_wire_412),
.PORT_ID_CLK(fresh_wire_411),
.PORT_ID_IN(fresh_wire_409),
.PORT_ID_OUT(fresh_wire_410));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(16'h0000),
.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3726$reg0(.PORT_ID_ARST(fresh_wire_416),
.PORT_ID_CLK(fresh_wire_415),
.PORT_ID_IN(fresh_wire_413),
.PORT_ID_OUT(fresh_wire_414));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(16'h0000),
.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3727$reg0(.PORT_ID_ARST(fresh_wire_420),
.PORT_ID_CLK(fresh_wire_419),
.PORT_ID_IN(fresh_wire_417),
.PORT_ID_OUT(fresh_wire_418));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3728$reg0(.PORT_ID_ARST(fresh_wire_424),
.PORT_ID_CLK(fresh_wire_423),
.PORT_ID_IN(fresh_wire_421),
.PORT_ID_OUT(fresh_wire_422));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3729$reg0(.PORT_ID_ARST(fresh_wire_428),
.PORT_ID_CLK(fresh_wire_427),
.PORT_ID_IN(fresh_wire_425),
.PORT_ID_OUT(fresh_wire_426));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3730$reg0(.PORT_ID_ARST(fresh_wire_432),
.PORT_ID_CLK(fresh_wire_431),
.PORT_ID_IN(fresh_wire_429),
.PORT_ID_OUT(fresh_wire_430));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2788$mux0(.PORT_ID_IN0(fresh_wire_433),
.PORT_ID_IN1(fresh_wire_434),
.PORT_ID_OUT(fresh_wire_435),
.PORT_ID_SEL(fresh_wire_436));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2865$mux0(.PORT_ID_IN0(fresh_wire_437),
.PORT_ID_IN1(fresh_wire_438),
.PORT_ID_OUT(fresh_wire_439),
.PORT_ID_SEL(fresh_wire_440));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2867$mux0(.PORT_ID_IN0(fresh_wire_441),
.PORT_ID_IN1(fresh_wire_442),
.PORT_ID_OUT(fresh_wire_443),
.PORT_ID_SEL(fresh_wire_444));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2877$mux0(.PORT_ID_IN0(fresh_wire_445),
.PORT_ID_IN1(fresh_wire_446),
.PORT_ID_OUT(fresh_wire_447),
.PORT_ID_SEL(fresh_wire_448));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2879$mux0(.PORT_ID_IN0(fresh_wire_449),
.PORT_ID_IN1(fresh_wire_450),
.PORT_ID_OUT(fresh_wire_451),
.PORT_ID_SEL(fresh_wire_452));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2888$mux0(.PORT_ID_IN0(fresh_wire_453),
.PORT_ID_IN1(fresh_wire_454),
.PORT_ID_OUT(fresh_wire_455),
.PORT_ID_SEL(fresh_wire_456));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2898$mux0(.PORT_ID_IN0(fresh_wire_457),
.PORT_ID_IN1(fresh_wire_458),
.PORT_ID_OUT(fresh_wire_459),
.PORT_ID_SEL(fresh_wire_460));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2904$mux0(.PORT_ID_IN0(fresh_wire_461),
.PORT_ID_IN1(fresh_wire_462),
.PORT_ID_OUT(fresh_wire_463),
.PORT_ID_SEL(fresh_wire_464));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2907$mux0(.PORT_ID_IN0(fresh_wire_465),
.PORT_ID_IN1(fresh_wire_466),
.PORT_ID_OUT(fresh_wire_467),
.PORT_ID_SEL(fresh_wire_468));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2909$mux0(.PORT_ID_IN0(fresh_wire_469),
.PORT_ID_IN1(fresh_wire_470),
.PORT_ID_OUT(fresh_wire_471),
.PORT_ID_SEL(fresh_wire_472));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2919$mux0(.PORT_ID_IN0(fresh_wire_473),
.PORT_ID_IN1(fresh_wire_474),
.PORT_ID_OUT(fresh_wire_475),
.PORT_ID_SEL(fresh_wire_476));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2923$mux0(.PORT_ID_IN0(fresh_wire_477),
.PORT_ID_IN1(fresh_wire_478),
.PORT_ID_OUT(fresh_wire_479),
.PORT_ID_SEL(fresh_wire_480));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2925$mux0(.PORT_ID_IN0(fresh_wire_481),
.PORT_ID_IN1(fresh_wire_482),
.PORT_ID_OUT(fresh_wire_483),
.PORT_ID_SEL(fresh_wire_484));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2931$mux0(.PORT_ID_IN0(fresh_wire_485),
.PORT_ID_IN1(fresh_wire_486),
.PORT_ID_OUT(fresh_wire_487),
.PORT_ID_SEL(fresh_wire_488));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2934$mux0(.PORT_ID_IN0(fresh_wire_489),
.PORT_ID_IN1(fresh_wire_490),
.PORT_ID_OUT(fresh_wire_491),
.PORT_ID_SEL(fresh_wire_492));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2936$mux0(.PORT_ID_IN0(fresh_wire_493),
.PORT_ID_IN1(fresh_wire_494),
.PORT_ID_OUT(fresh_wire_495),
.PORT_ID_SEL(fresh_wire_496));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2946$mux0(.PORT_ID_IN0(fresh_wire_497),
.PORT_ID_IN1(fresh_wire_498),
.PORT_ID_OUT(fresh_wire_499),
.PORT_ID_SEL(fresh_wire_500));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2952$mux0(.PORT_ID_IN0(fresh_wire_501),
.PORT_ID_IN1(fresh_wire_502),
.PORT_ID_OUT(fresh_wire_503),
.PORT_ID_SEL(fresh_wire_504));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2955$mux0(.PORT_ID_IN0(fresh_wire_505),
.PORT_ID_IN1(fresh_wire_506),
.PORT_ID_OUT(fresh_wire_507),
.PORT_ID_SEL(fresh_wire_508));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2957$mux0(.PORT_ID_IN0(fresh_wire_509),
.PORT_ID_IN1(fresh_wire_510),
.PORT_ID_OUT(fresh_wire_511),
.PORT_ID_SEL(fresh_wire_512));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2967$mux0(.PORT_ID_IN0(fresh_wire_513),
.PORT_ID_IN1(fresh_wire_514),
.PORT_ID_OUT(fresh_wire_515),
.PORT_ID_SEL(fresh_wire_516));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2971$mux0(.PORT_ID_IN0(fresh_wire_517),
.PORT_ID_IN1(fresh_wire_518),
.PORT_ID_OUT(fresh_wire_519),
.PORT_ID_SEL(fresh_wire_520));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2973$mux0(.PORT_ID_IN0(fresh_wire_521),
.PORT_ID_IN1(fresh_wire_522),
.PORT_ID_OUT(fresh_wire_523),
.PORT_ID_SEL(fresh_wire_524));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2979$mux0(.PORT_ID_IN0(fresh_wire_525),
.PORT_ID_IN1(fresh_wire_526),
.PORT_ID_OUT(fresh_wire_527),
.PORT_ID_SEL(fresh_wire_528));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2982$mux0(.PORT_ID_IN0(fresh_wire_529),
.PORT_ID_IN1(fresh_wire_530),
.PORT_ID_OUT(fresh_wire_531),
.PORT_ID_SEL(fresh_wire_532));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2984$mux0(.PORT_ID_IN0(fresh_wire_533),
.PORT_ID_IN1(fresh_wire_534),
.PORT_ID_OUT(fresh_wire_535),
.PORT_ID_SEL(fresh_wire_536));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2993$mux0(.PORT_ID_IN0(fresh_wire_537),
.PORT_ID_IN1(fresh_wire_538),
.PORT_ID_OUT(fresh_wire_539),
.PORT_ID_SEL(fresh_wire_540));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2997$mux0(.PORT_ID_IN0(fresh_wire_541),
.PORT_ID_IN1(fresh_wire_542),
.PORT_ID_OUT(fresh_wire_543),
.PORT_ID_SEL(fresh_wire_544));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2999$mux0(.PORT_ID_IN0(fresh_wire_545),
.PORT_ID_IN1(fresh_wire_546),
.PORT_ID_OUT(fresh_wire_547),
.PORT_ID_SEL(fresh_wire_548));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3013$mux0(.PORT_ID_IN0(fresh_wire_549),
.PORT_ID_IN1(fresh_wire_550),
.PORT_ID_OUT(fresh_wire_551),
.PORT_ID_SEL(fresh_wire_552));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3015$mux0(.PORT_ID_IN0(fresh_wire_553),
.PORT_ID_IN1(fresh_wire_554),
.PORT_ID_OUT(fresh_wire_555),
.PORT_ID_SEL(fresh_wire_556));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3017$mux0(.PORT_ID_IN0(fresh_wire_557),
.PORT_ID_IN1(fresh_wire_558),
.PORT_ID_OUT(fresh_wire_559),
.PORT_ID_SEL(fresh_wire_560));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3033$mux0(.PORT_ID_IN0(fresh_wire_561),
.PORT_ID_IN1(fresh_wire_562),
.PORT_ID_OUT(fresh_wire_563),
.PORT_ID_SEL(fresh_wire_564));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3035$mux0(.PORT_ID_IN0(fresh_wire_565),
.PORT_ID_IN1(fresh_wire_566),
.PORT_ID_OUT(fresh_wire_567),
.PORT_ID_SEL(fresh_wire_568));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3038$mux0(.PORT_ID_IN0(fresh_wire_569),
.PORT_ID_IN1(fresh_wire_570),
.PORT_ID_OUT(fresh_wire_571),
.PORT_ID_SEL(fresh_wire_572));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3057$mux0(.PORT_ID_IN0(fresh_wire_573),
.PORT_ID_IN1(fresh_wire_574),
.PORT_ID_OUT(fresh_wire_575),
.PORT_ID_SEL(fresh_wire_576));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3059$mux0(.PORT_ID_IN0(fresh_wire_577),
.PORT_ID_IN1(fresh_wire_578),
.PORT_ID_OUT(fresh_wire_579),
.PORT_ID_SEL(fresh_wire_580));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3069$mux0(.PORT_ID_IN0(fresh_wire_581),
.PORT_ID_IN1(fresh_wire_582),
.PORT_ID_OUT(fresh_wire_583),
.PORT_ID_SEL(fresh_wire_584));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3072$mux0(.PORT_ID_IN0(fresh_wire_585),
.PORT_ID_IN1(fresh_wire_586),
.PORT_ID_OUT(fresh_wire_587),
.PORT_ID_SEL(fresh_wire_588));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3074$mux0(.PORT_ID_IN0(fresh_wire_589),
.PORT_ID_IN1(fresh_wire_590),
.PORT_ID_OUT(fresh_wire_591),
.PORT_ID_SEL(fresh_wire_592));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__sub__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__244__DOLLAR__505$extendA(.PORT_ID_IN(fresh_wire_593),
.PORT_ID_OUT(fresh_wire_594));

	CELL_TYPE_SUB #(.PARAM_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__sub__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__244__DOLLAR__505$op0(.PORT_ID_IN0(fresh_wire_595),
.PORT_ID_IN1(fresh_wire_596),
.PORT_ID_OUT(fresh_wire_597));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__ternary__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__176__DOLLAR__475$mux0(.PORT_ID_IN0(fresh_wire_598),
.PORT_ID_IN1(fresh_wire_599),
.PORT_ID_OUT(fresh_wire_600),
.PORT_ID_SEL(fresh_wire_601));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__ternary__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__273__DOLLAR__526$mux0(.PORT_ID_IN0(fresh_wire_602),
.PORT_ID_IN1(fresh_wire_603),
.PORT_ID_OUT(fresh_wire_604),
.PORT_ID_SEL(fresh_wire_605));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__ternary__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__273__DOLLAR__526__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(.PORT_ID_OUT(fresh_wire_606));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$__DOLLAR__ternary__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__355__DOLLAR__569$mux0(.PORT_ID_IN0(fresh_wire_607),
.PORT_ID_IN1(fresh_wire_608),
.PORT_ID_OUT(fresh_wire_609),
.PORT_ID_SEL(fresh_wire_610));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__101__DOLLAR__314$op0(.PORT_ID_IN0(fresh_wire_611),
.PORT_ID_IN1(fresh_wire_612),
.PORT_ID_OUT(fresh_wire_613));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__100__DOLLAR__310$op0(.PORT_ID_IN0(fresh_wire_614),
.PORT_ID_IN1(fresh_wire_615),
.PORT_ID_OUT(fresh_wire_616));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__100__DOLLAR__311$op0(.PORT_ID_IN0(fresh_wire_617),
.PORT_ID_IN1(fresh_wire_618),
.PORT_ID_OUT(fresh_wire_619));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__103__DOLLAR__316$op0(.PORT_ID_IN0(fresh_wire_620),
.PORT_ID_IN1(fresh_wire_621),
.PORT_ID_OUT(fresh_wire_622));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__128__DOLLAR__345$op0(.PORT_ID_IN0(fresh_wire_623),
.PORT_ID_IN1(fresh_wire_624),
.PORT_ID_OUT(fresh_wire_625));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__150__DOLLAR__379$op0(.PORT_ID_IN0(fresh_wire_626),
.PORT_ID_IN1(fresh_wire_627),
.PORT_ID_OUT(fresh_wire_628));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__157__DOLLAR__381$op0(.PORT_ID_IN0(fresh_wire_629),
.PORT_ID_IN1(fresh_wire_630),
.PORT_ID_OUT(fresh_wire_631));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__158__DOLLAR__382$op0(.PORT_ID_IN0(fresh_wire_632),
.PORT_ID_IN1(fresh_wire_633),
.PORT_ID_OUT(fresh_wire_634));

	CELL_TYPE_UGE #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__ge__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__126__DOLLAR__341$op0(.PORT_ID_IN0(fresh_wire_635),
.PORT_ID_IN1(fresh_wire_636),
.PORT_ID_OUT(fresh_wire_637));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__100__DOLLAR__312$aRed(.PORT_ID_IN(fresh_wire_638),
.PORT_ID_OUT(fresh_wire_639));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__100__DOLLAR__312$andOps(.PORT_ID_IN0(fresh_wire_640),
.PORT_ID_IN1(fresh_wire_641),
.PORT_ID_OUT(fresh_wire_642));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__100__DOLLAR__312$bRed(.PORT_ID_IN(fresh_wire_643),
.PORT_ID_OUT(fresh_wire_644));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__100__DOLLAR__313$andOps(.PORT_ID_IN0(fresh_wire_645),
.PORT_ID_IN1(fresh_wire_646),
.PORT_ID_OUT(fresh_wire_647));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__100__DOLLAR__313$bRed(.PORT_ID_IN(fresh_wire_648),
.PORT_ID_OUT(fresh_wire_649));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__103__DOLLAR__317$andOps(.PORT_ID_IN0(fresh_wire_650),
.PORT_ID_IN1(fresh_wire_651),
.PORT_ID_OUT(fresh_wire_652));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__103__DOLLAR__317$bRed(.PORT_ID_IN(fresh_wire_653),
.PORT_ID_OUT(fresh_wire_654));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__125__DOLLAR__340$andOps(.PORT_ID_IN0(fresh_wire_655),
.PORT_ID_IN1(fresh_wire_656),
.PORT_ID_OUT(fresh_wire_657));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__125__DOLLAR__340$bRed(.PORT_ID_IN(fresh_wire_658),
.PORT_ID_OUT(fresh_wire_659));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__127__DOLLAR__344$andOps(.PORT_ID_IN0(fresh_wire_660),
.PORT_ID_IN1(fresh_wire_661),
.PORT_ID_OUT(fresh_wire_662));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__127__DOLLAR__344$bRed(.PORT_ID_IN(fresh_wire_663),
.PORT_ID_OUT(fresh_wire_664));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(2'h0),
.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__procdff__DOLLAR__3739$reg0(.PORT_ID_ARST(fresh_wire_668),
.PORT_ID_CLK(fresh_wire_667),
.PORT_ID_IN(fresh_wire_665),
.PORT_ID_OUT(fresh_wire_666));

	CELL_TYPE_REG #(.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(48'hxxxxxxxxxxxx),
.PARAM_WIDTH(32'h00000030)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__procdff__DOLLAR__3740$reg0(.PORT_ID_CLK(fresh_wire_671),
.PORT_ID_IN(fresh_wire_669),
.PORT_ID_OUT(fresh_wire_670));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3178$mux0(.PORT_ID_IN0(fresh_wire_672),
.PORT_ID_IN1(fresh_wire_673),
.PORT_ID_OUT(fresh_wire_674),
.PORT_ID_SEL(fresh_wire_675));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3181$mux0(.PORT_ID_IN0(fresh_wire_676),
.PORT_ID_IN1(fresh_wire_677),
.PORT_ID_OUT(fresh_wire_678),
.PORT_ID_SEL(fresh_wire_679));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3199$mux0(.PORT_ID_IN0(fresh_wire_680),
.PORT_ID_IN1(fresh_wire_681),
.PORT_ID_OUT(fresh_wire_682),
.PORT_ID_SEL(fresh_wire_683));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3202$mux0(.PORT_ID_IN0(fresh_wire_684),
.PORT_ID_IN1(fresh_wire_685),
.PORT_ID_OUT(fresh_wire_686),
.PORT_ID_SEL(fresh_wire_687));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3211$mux0(.PORT_ID_IN0(fresh_wire_688),
.PORT_ID_IN1(fresh_wire_689),
.PORT_ID_OUT(fresh_wire_690),
.PORT_ID_SEL(fresh_wire_691));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3214$mux0(.PORT_ID_IN0(fresh_wire_692),
.PORT_ID_IN1(fresh_wire_693),
.PORT_ID_OUT(fresh_wire_694),
.PORT_ID_SEL(fresh_wire_695));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3217$mux0(.PORT_ID_IN0(fresh_wire_696),
.PORT_ID_IN1(fresh_wire_697),
.PORT_ID_OUT(fresh_wire_698),
.PORT_ID_SEL(fresh_wire_699));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3219$mux0(.PORT_ID_IN0(fresh_wire_700),
.PORT_ID_IN1(fresh_wire_701),
.PORT_ID_OUT(fresh_wire_702),
.PORT_ID_SEL(fresh_wire_703));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3223$mux0(.PORT_ID_IN0(fresh_wire_704),
.PORT_ID_IN1(fresh_wire_705),
.PORT_ID_OUT(fresh_wire_706),
.PORT_ID_SEL(fresh_wire_707));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3226$mux0(.PORT_ID_IN0(fresh_wire_708),
.PORT_ID_IN1(fresh_wire_709),
.PORT_ID_OUT(fresh_wire_710),
.PORT_ID_SEL(fresh_wire_711));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000020)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3228$mux0(.PORT_ID_IN0(fresh_wire_712),
.PORT_ID_IN1(fresh_wire_713),
.PORT_ID_OUT(fresh_wire_714),
.PORT_ID_SEL(fresh_wire_715));

	CELL_TYPE_SUB #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__sub__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__104__DOLLAR__318$op0(.PORT_ID_IN0(fresh_wire_716),
.PORT_ID_IN1(fresh_wire_717),
.PORT_ID_OUT(fresh_wire_718));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$input_sr$__DOLLAR__sub__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__110__DOLLAR__326__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(.PORT_ID_OUT(fresh_wire_719));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__103__DOLLAR__747$op0(.PORT_ID_IN0(fresh_wire_720),
.PORT_ID_IN1(fresh_wire_721),
.PORT_ID_OUT(fresh_wire_722));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__106__DOLLAR__751$op0(.PORT_ID_IN0(fresh_wire_723),
.PORT_ID_IN1(fresh_wire_724),
.PORT_ID_OUT(fresh_wire_725));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__102__DOLLAR__744$op0(.PORT_ID_IN0(fresh_wire_726),
.PORT_ID_IN1(fresh_wire_727),
.PORT_ID_OUT(fresh_wire_728));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__102__DOLLAR__745$op0(.PORT_ID_IN0(fresh_wire_729),
.PORT_ID_IN1(fresh_wire_730),
.PORT_ID_OUT(fresh_wire_731));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__105__DOLLAR__748$op0(.PORT_ID_IN0(fresh_wire_732),
.PORT_ID_IN1(fresh_wire_733),
.PORT_ID_OUT(fresh_wire_734));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__108__DOLLAR__753$op0(.PORT_ID_IN0(fresh_wire_735),
.PORT_ID_IN1(fresh_wire_736),
.PORT_ID_OUT(fresh_wire_737));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__120__DOLLAR__760$op0(.PORT_ID_IN0(fresh_wire_738),
.PORT_ID_IN1(fresh_wire_739),
.PORT_ID_OUT(fresh_wire_740));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__120__DOLLAR__761$op0(.PORT_ID_IN0(fresh_wire_741),
.PORT_ID_IN1(fresh_wire_742),
.PORT_ID_OUT(fresh_wire_743));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__133__DOLLAR__784$op0(.PORT_ID_IN0(fresh_wire_744),
.PORT_ID_IN1(fresh_wire_745),
.PORT_ID_OUT(fresh_wire_746));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__135__DOLLAR__785$op0(.PORT_ID_IN0(fresh_wire_747),
.PORT_ID_IN1(fresh_wire_748),
.PORT_ID_OUT(fresh_wire_749));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__137__DOLLAR__786$op0(.PORT_ID_IN0(fresh_wire_750),
.PORT_ID_IN1(fresh_wire_751),
.PORT_ID_OUT(fresh_wire_752));

	CELL_TYPE_UGE #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__ge__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__121__DOLLAR__765$op0(.PORT_ID_IN0(fresh_wire_753),
.PORT_ID_IN1(fresh_wire_754),
.PORT_ID_OUT(fresh_wire_755));

	CELL_TYPE_UGE #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__ge__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__123__DOLLAR__771$op0(.PORT_ID_IN0(fresh_wire_756),
.PORT_ID_IN1(fresh_wire_757),
.PORT_ID_OUT(fresh_wire_758));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__102__DOLLAR__746$aRed(.PORT_ID_IN(fresh_wire_759),
.PORT_ID_OUT(fresh_wire_760));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__102__DOLLAR__746$andOps(.PORT_ID_IN0(fresh_wire_761),
.PORT_ID_IN1(fresh_wire_762),
.PORT_ID_OUT(fresh_wire_763));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__102__DOLLAR__746$bRed(.PORT_ID_IN(fresh_wire_764),
.PORT_ID_OUT(fresh_wire_765));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__105__DOLLAR__750$aRed(.PORT_ID_IN(fresh_wire_766),
.PORT_ID_OUT(fresh_wire_767));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__105__DOLLAR__750$andOps(.PORT_ID_IN0(fresh_wire_768),
.PORT_ID_IN1(fresh_wire_769),
.PORT_ID_OUT(fresh_wire_770));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__105__DOLLAR__750$bRed(.PORT_ID_IN(fresh_wire_771),
.PORT_ID_OUT(fresh_wire_772));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__108__DOLLAR__754$aRed(.PORT_ID_IN(fresh_wire_773),
.PORT_ID_OUT(fresh_wire_774));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__108__DOLLAR__754$andOps(.PORT_ID_IN0(fresh_wire_775),
.PORT_ID_IN1(fresh_wire_776),
.PORT_ID_OUT(fresh_wire_777));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__108__DOLLAR__754$bRed(.PORT_ID_IN(fresh_wire_778),
.PORT_ID_OUT(fresh_wire_779));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__110__DOLLAR__757$aRed(.PORT_ID_IN(fresh_wire_780),
.PORT_ID_OUT(fresh_wire_781));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__110__DOLLAR__757$andOps(.PORT_ID_IN0(fresh_wire_782),
.PORT_ID_IN1(fresh_wire_783),
.PORT_ID_OUT(fresh_wire_784));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__110__DOLLAR__757$bRed(.PORT_ID_IN(fresh_wire_785),
.PORT_ID_OUT(fresh_wire_786));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__120__DOLLAR__762$aRed(.PORT_ID_IN(fresh_wire_787),
.PORT_ID_OUT(fresh_wire_788));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__120__DOLLAR__762$andOps(.PORT_ID_IN0(fresh_wire_789),
.PORT_ID_IN1(fresh_wire_790),
.PORT_ID_OUT(fresh_wire_791));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__120__DOLLAR__762$bRed(.PORT_ID_IN(fresh_wire_792),
.PORT_ID_OUT(fresh_wire_793));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__120__DOLLAR__764$aRed(.PORT_ID_IN(fresh_wire_794),
.PORT_ID_OUT(fresh_wire_795));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__120__DOLLAR__764$andOps(.PORT_ID_IN0(fresh_wire_796),
.PORT_ID_IN1(fresh_wire_797),
.PORT_ID_OUT(fresh_wire_798));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__120__DOLLAR__764$bRed(.PORT_ID_IN(fresh_wire_799),
.PORT_ID_OUT(fresh_wire_800));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__122__DOLLAR__768$aRed(.PORT_ID_IN(fresh_wire_801),
.PORT_ID_OUT(fresh_wire_802));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__122__DOLLAR__768$andOps(.PORT_ID_IN0(fresh_wire_803),
.PORT_ID_IN1(fresh_wire_804),
.PORT_ID_OUT(fresh_wire_805));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__122__DOLLAR__768$bRed(.PORT_ID_IN(fresh_wire_806),
.PORT_ID_OUT(fresh_wire_807));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__122__DOLLAR__770$aRed(.PORT_ID_IN(fresh_wire_808),
.PORT_ID_OUT(fresh_wire_809));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__122__DOLLAR__770$andOps(.PORT_ID_IN0(fresh_wire_810),
.PORT_ID_IN1(fresh_wire_811),
.PORT_ID_OUT(fresh_wire_812));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__122__DOLLAR__770$bRed(.PORT_ID_IN(fresh_wire_813),
.PORT_ID_OUT(fresh_wire_814));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__124__DOLLAR__776$aRed(.PORT_ID_IN(fresh_wire_815),
.PORT_ID_OUT(fresh_wire_816));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__124__DOLLAR__776$andOps(.PORT_ID_IN0(fresh_wire_817),
.PORT_ID_IN1(fresh_wire_818),
.PORT_ID_OUT(fresh_wire_819));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__124__DOLLAR__776$bRed(.PORT_ID_IN(fresh_wire_820),
.PORT_ID_OUT(fresh_wire_821));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__126__DOLLAR__781$aRed(.PORT_ID_IN(fresh_wire_822),
.PORT_ID_OUT(fresh_wire_823));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__126__DOLLAR__781$andOps(.PORT_ID_IN0(fresh_wire_824),
.PORT_ID_IN1(fresh_wire_825),
.PORT_ID_OUT(fresh_wire_826));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__126__DOLLAR__781$bRed(.PORT_ID_IN(fresh_wire_827),
.PORT_ID_OUT(fresh_wire_828));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__99__DOLLAR__740$aRed(.PORT_ID_IN(fresh_wire_829),
.PORT_ID_OUT(fresh_wire_830));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__99__DOLLAR__740$andOps(.PORT_ID_IN0(fresh_wire_831),
.PORT_ID_IN1(fresh_wire_832),
.PORT_ID_OUT(fresh_wire_833));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__99__DOLLAR__740$bRed(.PORT_ID_IN(fresh_wire_834),
.PORT_ID_OUT(fresh_wire_835));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__99__DOLLAR__742$aRed(.PORT_ID_IN(fresh_wire_836),
.PORT_ID_OUT(fresh_wire_837));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__99__DOLLAR__742$andOps(.PORT_ID_IN0(fresh_wire_838),
.PORT_ID_IN1(fresh_wire_839),
.PORT_ID_OUT(fresh_wire_840));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__99__DOLLAR__742$bRed(.PORT_ID_IN(fresh_wire_841),
.PORT_ID_OUT(fresh_wire_842));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_or__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__124__DOLLAR__774$aRed(.PORT_ID_IN(fresh_wire_843),
.PORT_ID_OUT(fresh_wire_844));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_or__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__124__DOLLAR__774$bRed(.PORT_ID_IN(fresh_wire_845),
.PORT_ID_OUT(fresh_wire_846));

	CELL_TYPE_OR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_or__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__124__DOLLAR__774$orOps(.PORT_ID_IN0(fresh_wire_847),
.PORT_ID_IN1(fresh_wire_848),
.PORT_ID_OUT(fresh_wire_849));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_or__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__126__DOLLAR__779$aRed(.PORT_ID_IN(fresh_wire_850),
.PORT_ID_OUT(fresh_wire_851));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_or__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__126__DOLLAR__779$bRed(.PORT_ID_IN(fresh_wire_852),
.PORT_ID_OUT(fresh_wire_853));

	CELL_TYPE_OR #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_or__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__126__DOLLAR__779$orOps(.PORT_ID_IN0(fresh_wire_854),
.PORT_ID_IN1(fresh_wire_855),
.PORT_ID_OUT(fresh_wire_856));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(2'h0),
.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procdff__DOLLAR__3701$reg0(.PORT_ID_ARST(fresh_wire_860),
.PORT_ID_CLK(fresh_wire_859),
.PORT_ID_IN(fresh_wire_857),
.PORT_ID_OUT(fresh_wire_858));

	CELL_TYPE_REG #(.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(48'hxxxxxxxxxxxx),
.PARAM_WIDTH(32'h00000030)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procdff__DOLLAR__3702$reg0(.PORT_ID_CLK(fresh_wire_863),
.PORT_ID_IN(fresh_wire_861),
.PORT_ID_OUT(fresh_wire_862));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2382$mux0(.PORT_ID_IN0(fresh_wire_864),
.PORT_ID_IN1(fresh_wire_865),
.PORT_ID_OUT(fresh_wire_866),
.PORT_ID_SEL(fresh_wire_867));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2385$mux0(.PORT_ID_IN0(fresh_wire_868),
.PORT_ID_IN1(fresh_wire_869),
.PORT_ID_OUT(fresh_wire_870),
.PORT_ID_SEL(fresh_wire_871));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2388$mux0(.PORT_ID_IN0(fresh_wire_872),
.PORT_ID_IN1(fresh_wire_873),
.PORT_ID_OUT(fresh_wire_874),
.PORT_ID_SEL(fresh_wire_875));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2390$mux0(.PORT_ID_IN0(fresh_wire_876),
.PORT_ID_IN1(fresh_wire_877),
.PORT_ID_OUT(fresh_wire_878),
.PORT_ID_SEL(fresh_wire_879));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2393$mux0(.PORT_ID_IN0(fresh_wire_880),
.PORT_ID_IN1(fresh_wire_881),
.PORT_ID_OUT(fresh_wire_882),
.PORT_ID_SEL(fresh_wire_883));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2396$mux0(.PORT_ID_IN0(fresh_wire_884),
.PORT_ID_IN1(fresh_wire_885),
.PORT_ID_OUT(fresh_wire_886),
.PORT_ID_SEL(fresh_wire_887));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2399$mux0(.PORT_ID_IN0(fresh_wire_888),
.PORT_ID_IN1(fresh_wire_889),
.PORT_ID_OUT(fresh_wire_890),
.PORT_ID_SEL(fresh_wire_891));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2402$mux0(.PORT_ID_IN0(fresh_wire_892),
.PORT_ID_IN1(fresh_wire_893),
.PORT_ID_OUT(fresh_wire_894),
.PORT_ID_SEL(fresh_wire_895));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2406$mux0(.PORT_ID_IN0(fresh_wire_896),
.PORT_ID_IN1(fresh_wire_897),
.PORT_ID_OUT(fresh_wire_898),
.PORT_ID_SEL(fresh_wire_899));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2409$mux0(.PORT_ID_IN0(fresh_wire_900),
.PORT_ID_IN1(fresh_wire_901),
.PORT_ID_OUT(fresh_wire_902),
.PORT_ID_SEL(fresh_wire_903));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2412$mux0(.PORT_ID_IN0(fresh_wire_904),
.PORT_ID_IN1(fresh_wire_905),
.PORT_ID_OUT(fresh_wire_906),
.PORT_ID_SEL(fresh_wire_907));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2415$mux0(.PORT_ID_IN0(fresh_wire_908),
.PORT_ID_IN1(fresh_wire_909),
.PORT_ID_OUT(fresh_wire_910),
.PORT_ID_SEL(fresh_wire_911));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2418$mux0(.PORT_ID_IN0(fresh_wire_912),
.PORT_ID_IN1(fresh_wire_913),
.PORT_ID_OUT(fresh_wire_914),
.PORT_ID_SEL(fresh_wire_915));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000030)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2427$mux0(.PORT_ID_IN0(fresh_wire_916),
.PORT_ID_IN1(fresh_wire_917),
.PORT_ID_OUT(fresh_wire_918),
.PORT_ID_SEL(fresh_wire_919));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000030)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2430$mux0(.PORT_ID_IN0(fresh_wire_920),
.PORT_ID_IN1(fresh_wire_921),
.PORT_ID_OUT(fresh_wire_922),
.PORT_ID_SEL(fresh_wire_923));

	CELL_TYPE_SUB #(.PARAM_WIDTH(32'h00000002)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__sub__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__100__DOLLAR__743$op0(.PORT_ID_IN0(fresh_wire_924),
.PORT_ID_IN1(fresh_wire_925),
.PORT_ID_OUT(fresh_wire_926));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$linebuffer_control$output_sr$__DOLLAR__sub__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__100__DOLLAR__743__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(.PORT_ID_OUT(fresh_wire_927));

	CELL_TYPE_NOT #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$__DOLLAR__not__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__mem_unq1__DOT__v__COLON__65__DOLLAR__575$op0(.PORT_ID_IN(fresh_wire_928),
.PORT_ID_OUT(fresh_wire_929));

	CELL_TYPE_NOT #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$__DOLLAR__not__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__mem_unq1__DOT__v__COLON__66__DOLLAR__576$op0(.PORT_ID_IN(fresh_wire_930),
.PORT_ID_OUT(fresh_wire_931));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__sram_512w_16b__DOT__v__COLON__38__DOLLAR__1114$op0(.PORT_ID_IN0(fresh_wire_932),
.PORT_ID_IN1(fresh_wire_933),
.PORT_ID_OUT(fresh_wire_934));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__sram_512w_16b__DOT__v__COLON__40__DOLLAR__1116$op0(.PORT_ID_IN0(fresh_wire_935),
.PORT_ID_IN1(fresh_wire_936),
.PORT_ID_OUT(fresh_wire_937));

	CELL_TYPE_REG #(.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(16'hxxxx),
.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procdff__DOLLAR__3630$reg0(.PORT_ID_CLK(fresh_wire_940),
.PORT_ID_IN(fresh_wire_938),
.PORT_ID_OUT(fresh_wire_939));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1557$mux0(.PORT_ID_IN0(fresh_wire_941),
.PORT_ID_IN1(fresh_wire_942),
.PORT_ID_OUT(fresh_wire_943),
.PORT_ID_SEL(fresh_wire_944));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1567$mux0(.PORT_ID_IN0(fresh_wire_945),
.PORT_ID_IN1(fresh_wire_946),
.PORT_ID_OUT(fresh_wire_947),
.PORT_ID_SEL(fresh_wire_948));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1567__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(.PORT_ID_OUT(fresh_wire_949));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1569$mux0(.PORT_ID_IN0(fresh_wire_950),
.PORT_ID_IN1(fresh_wire_951),
.PORT_ID_OUT(fresh_wire_952),
.PORT_ID_SEL(fresh_wire_953));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576$mux0(.PORT_ID_IN0(fresh_wire_954),
.PORT_ID_IN1(fresh_wire_955),
.PORT_ID_OUT(fresh_wire_956),
.PORT_ID_SEL(fresh_wire_957));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0$uConst(.PORT_ID_OUT(fresh_wire_958));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10$uConst(.PORT_ID_OUT(fresh_wire_959));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11$uConst(.PORT_ID_OUT(fresh_wire_960));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12$uConst(.PORT_ID_OUT(fresh_wire_961));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13$uConst(.PORT_ID_OUT(fresh_wire_962));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14$uConst(.PORT_ID_OUT(fresh_wire_963));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15$uConst(.PORT_ID_OUT(fresh_wire_964));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1$uConst(.PORT_ID_OUT(fresh_wire_965));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2$uConst(.PORT_ID_OUT(fresh_wire_966));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3$uConst(.PORT_ID_OUT(fresh_wire_967));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4$uConst(.PORT_ID_OUT(fresh_wire_968));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5$uConst(.PORT_ID_OUT(fresh_wire_969));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6$uConst(.PORT_ID_OUT(fresh_wire_970));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7$uConst(.PORT_ID_OUT(fresh_wire_971));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8$uConst(.PORT_ID_OUT(fresh_wire_972));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9$uConst(.PORT_ID_OUT(fresh_wire_973));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578$mux0(.PORT_ID_IN0(fresh_wire_974),
.PORT_ID_IN1(fresh_wire_975),
.PORT_ID_OUT(fresh_wire_976),
.PORT_ID_SEL(fresh_wire_977));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0$uConst(.PORT_ID_OUT(fresh_wire_978));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10$uConst(.PORT_ID_OUT(fresh_wire_979));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11$uConst(.PORT_ID_OUT(fresh_wire_980));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12$uConst(.PORT_ID_OUT(fresh_wire_981));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13$uConst(.PORT_ID_OUT(fresh_wire_982));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14$uConst(.PORT_ID_OUT(fresh_wire_983));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15$uConst(.PORT_ID_OUT(fresh_wire_984));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1$uConst(.PORT_ID_OUT(fresh_wire_985));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2$uConst(.PORT_ID_OUT(fresh_wire_986));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3$uConst(.PORT_ID_OUT(fresh_wire_987));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4$uConst(.PORT_ID_OUT(fresh_wire_988));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5$uConst(.PORT_ID_OUT(fresh_wire_989));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6$uConst(.PORT_ID_OUT(fresh_wire_990));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7$uConst(.PORT_ID_OUT(fresh_wire_991));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8$uConst(.PORT_ID_OUT(fresh_wire_992));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9$uConst(.PORT_ID_OUT(fresh_wire_993));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000009)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585$mux0(.PORT_ID_IN0(fresh_wire_994),
.PORT_ID_IN1(fresh_wire_995),
.PORT_ID_OUT(fresh_wire_996),
.PORT_ID_SEL(fresh_wire_997));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0$uConst(.PORT_ID_OUT(fresh_wire_998));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1$uConst(.PORT_ID_OUT(fresh_wire_999));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2$uConst(.PORT_ID_OUT(fresh_wire_1000));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3$uConst(.PORT_ID_OUT(fresh_wire_1001));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4$uConst(.PORT_ID_OUT(fresh_wire_1002));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5$uConst(.PORT_ID_OUT(fresh_wire_1003));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6$uConst(.PORT_ID_OUT(fresh_wire_1004));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7$uConst(.PORT_ID_OUT(fresh_wire_1005));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8$uConst(.PORT_ID_OUT(fresh_wire_1006));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000009)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587$mux0(.PORT_ID_IN0(fresh_wire_1007),
.PORT_ID_IN1(fresh_wire_1008),
.PORT_ID_OUT(fresh_wire_1009),
.PORT_ID_SEL(fresh_wire_1010));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0$uConst(.PORT_ID_OUT(fresh_wire_1011));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1$uConst(.PORT_ID_OUT(fresh_wire_1012));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2$uConst(.PORT_ID_OUT(fresh_wire_1013));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3$uConst(.PORT_ID_OUT(fresh_wire_1014));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4$uConst(.PORT_ID_OUT(fresh_wire_1015));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5$uConst(.PORT_ID_OUT(fresh_wire_1016));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6$uConst(.PORT_ID_OUT(fresh_wire_1017));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7$uConst(.PORT_ID_OUT(fresh_wire_1018));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8$uConst(.PORT_ID_OUT(fresh_wire_1019));

	CELL_TYPE_MEM #(.PARAM_HAS_INIT(1'h0),
.PARAM_MEM_DEPTH(32'h00000200),
.PARAM_MEM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst0$mem_inst$data_array$mem(.PORT_ID_CLK(fresh_wire_1020),
.PORT_ID_RADDR(fresh_wire_1021),
.PORT_ID_RDATA(fresh_wire_1022),
.PORT_ID_WADDR(fresh_wire_1023),
.PORT_ID_WDATA(fresh_wire_1024),
.PORT_ID_WEN(fresh_wire_1025));

	CELL_TYPE_NOT #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$__DOLLAR__not__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__mem_unq1__DOT__v__COLON__65__DOLLAR__575$op0(.PORT_ID_IN(fresh_wire_1026),
.PORT_ID_OUT(fresh_wire_1027));

	CELL_TYPE_NOT #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$__DOLLAR__not__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__mem_unq1__DOT__v__COLON__66__DOLLAR__576$op0(.PORT_ID_IN(fresh_wire_1028),
.PORT_ID_OUT(fresh_wire_1029));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__sram_512w_16b__DOT__v__COLON__38__DOLLAR__1114$op0(.PORT_ID_IN0(fresh_wire_1030),
.PORT_ID_IN1(fresh_wire_1031),
.PORT_ID_OUT(fresh_wire_1032));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__sram_512w_16b__DOT__v__COLON__40__DOLLAR__1116$op0(.PORT_ID_IN0(fresh_wire_1033),
.PORT_ID_IN1(fresh_wire_1034),
.PORT_ID_OUT(fresh_wire_1035));

	CELL_TYPE_REG #(.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(16'hxxxx),
.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procdff__DOLLAR__3630$reg0(.PORT_ID_CLK(fresh_wire_1038),
.PORT_ID_IN(fresh_wire_1036),
.PORT_ID_OUT(fresh_wire_1037));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1557$mux0(.PORT_ID_IN0(fresh_wire_1039),
.PORT_ID_IN1(fresh_wire_1040),
.PORT_ID_OUT(fresh_wire_1041),
.PORT_ID_SEL(fresh_wire_1042));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1567$mux0(.PORT_ID_IN0(fresh_wire_1043),
.PORT_ID_IN1(fresh_wire_1044),
.PORT_ID_OUT(fresh_wire_1045),
.PORT_ID_SEL(fresh_wire_1046));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1567__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(.PORT_ID_OUT(fresh_wire_1047));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1569$mux0(.PORT_ID_IN0(fresh_wire_1048),
.PORT_ID_IN1(fresh_wire_1049),
.PORT_ID_OUT(fresh_wire_1050),
.PORT_ID_SEL(fresh_wire_1051));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576$mux0(.PORT_ID_IN0(fresh_wire_1052),
.PORT_ID_IN1(fresh_wire_1053),
.PORT_ID_OUT(fresh_wire_1054),
.PORT_ID_SEL(fresh_wire_1055));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0$uConst(.PORT_ID_OUT(fresh_wire_1056));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10$uConst(.PORT_ID_OUT(fresh_wire_1057));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11$uConst(.PORT_ID_OUT(fresh_wire_1058));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12$uConst(.PORT_ID_OUT(fresh_wire_1059));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13$uConst(.PORT_ID_OUT(fresh_wire_1060));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14$uConst(.PORT_ID_OUT(fresh_wire_1061));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15$uConst(.PORT_ID_OUT(fresh_wire_1062));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1$uConst(.PORT_ID_OUT(fresh_wire_1063));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2$uConst(.PORT_ID_OUT(fresh_wire_1064));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3$uConst(.PORT_ID_OUT(fresh_wire_1065));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4$uConst(.PORT_ID_OUT(fresh_wire_1066));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5$uConst(.PORT_ID_OUT(fresh_wire_1067));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6$uConst(.PORT_ID_OUT(fresh_wire_1068));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7$uConst(.PORT_ID_OUT(fresh_wire_1069));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8$uConst(.PORT_ID_OUT(fresh_wire_1070));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9$uConst(.PORT_ID_OUT(fresh_wire_1071));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578$mux0(.PORT_ID_IN0(fresh_wire_1072),
.PORT_ID_IN1(fresh_wire_1073),
.PORT_ID_OUT(fresh_wire_1074),
.PORT_ID_SEL(fresh_wire_1075));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0$uConst(.PORT_ID_OUT(fresh_wire_1076));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10$uConst(.PORT_ID_OUT(fresh_wire_1077));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11$uConst(.PORT_ID_OUT(fresh_wire_1078));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12$uConst(.PORT_ID_OUT(fresh_wire_1079));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13$uConst(.PORT_ID_OUT(fresh_wire_1080));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14$uConst(.PORT_ID_OUT(fresh_wire_1081));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15$uConst(.PORT_ID_OUT(fresh_wire_1082));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1$uConst(.PORT_ID_OUT(fresh_wire_1083));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2$uConst(.PORT_ID_OUT(fresh_wire_1084));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3$uConst(.PORT_ID_OUT(fresh_wire_1085));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4$uConst(.PORT_ID_OUT(fresh_wire_1086));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5$uConst(.PORT_ID_OUT(fresh_wire_1087));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6$uConst(.PORT_ID_OUT(fresh_wire_1088));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7$uConst(.PORT_ID_OUT(fresh_wire_1089));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8$uConst(.PORT_ID_OUT(fresh_wire_1090));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9$uConst(.PORT_ID_OUT(fresh_wire_1091));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000009)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585$mux0(.PORT_ID_IN0(fresh_wire_1092),
.PORT_ID_IN1(fresh_wire_1093),
.PORT_ID_OUT(fresh_wire_1094),
.PORT_ID_SEL(fresh_wire_1095));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0$uConst(.PORT_ID_OUT(fresh_wire_1096));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1$uConst(.PORT_ID_OUT(fresh_wire_1097));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2$uConst(.PORT_ID_OUT(fresh_wire_1098));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3$uConst(.PORT_ID_OUT(fresh_wire_1099));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4$uConst(.PORT_ID_OUT(fresh_wire_1100));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5$uConst(.PORT_ID_OUT(fresh_wire_1101));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6$uConst(.PORT_ID_OUT(fresh_wire_1102));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7$uConst(.PORT_ID_OUT(fresh_wire_1103));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8$uConst(.PORT_ID_OUT(fresh_wire_1104));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000009)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587$mux0(.PORT_ID_IN0(fresh_wire_1105),
.PORT_ID_IN1(fresh_wire_1106),
.PORT_ID_OUT(fresh_wire_1107),
.PORT_ID_SEL(fresh_wire_1108));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0$uConst(.PORT_ID_OUT(fresh_wire_1109));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1$uConst(.PORT_ID_OUT(fresh_wire_1110));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2$uConst(.PORT_ID_OUT(fresh_wire_1111));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3$uConst(.PORT_ID_OUT(fresh_wire_1112));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4$uConst(.PORT_ID_OUT(fresh_wire_1113));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5$uConst(.PORT_ID_OUT(fresh_wire_1114));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6$uConst(.PORT_ID_OUT(fresh_wire_1115));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7$uConst(.PORT_ID_OUT(fresh_wire_1116));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x18$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8$uConst(.PORT_ID_OUT(fresh_wire_1117));

	CELL_TYPE_MEM #(.PARAM_HAS_INIT(1'h0),
.PARAM_MEM_DEPTH(32'h00000200),
.PARAM_MEM_WIDTH(32'h00000010)) mem_0x18$memory_core$mem_inst1$mem_inst$data_array$mem(.PORT_ID_CLK(fresh_wire_1118),
.PORT_ID_RADDR(fresh_wire_1119),
.PORT_ID_RDATA(fresh_wire_1120),
.PORT_ID_WADDR(fresh_wire_1121),
.PORT_ID_WDATA(fresh_wire_1122),
.PORT_ID_WEN(fresh_wire_1123));

	CELL_TYPE_REG #(.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(16'hxxxx),
.PARAM_WIDTH(32'h00000010)) mem_0x18$sb_inst_busBUS16_row0$__DOLLAR__procdff__DOLLAR__3697$reg0(.PORT_ID_CLK(fresh_wire_1126),
.PORT_ID_IN(fresh_wire_1124),
.PORT_ID_OUT(fresh_wire_1125));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$__DOLLAR__and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__memory_core_unq1__DOT__v__COLON__309__DOLLAR__631$op0(.PORT_ID_IN0(fresh_wire_1127),
.PORT_ID_IN1(fresh_wire_1128),
.PORT_ID_OUT(fresh_wire_1129));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$__DOLLAR__and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__memory_core_unq1__DOT__v__COLON__310__DOLLAR__633$op0(.PORT_ID_IN0(fresh_wire_1130),
.PORT_ID_IN1(fresh_wire_1131),
.PORT_ID_OUT(fresh_wire_1132));

	CELL_TYPE_OR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$__DOLLAR__or__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__memory_core_unq1__DOT__v__COLON__309__DOLLAR__630$op0(.PORT_ID_IN0(fresh_wire_1133),
.PORT_ID_IN1(fresh_wire_1134),
.PORT_ID_OUT(fresh_wire_1135));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__471$op0(.PORT_ID_IN0(fresh_wire_1136),
.PORT_ID_IN1(fresh_wire_1137),
.PORT_ID_OUT(fresh_wire_1138));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000002),
.PARAM_OUT_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__206__DOLLAR__488$extendB(.PORT_ID_IN(fresh_wire_1139),
.PORT_ID_OUT(fresh_wire_1140));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__206__DOLLAR__488$op0(.PORT_ID_IN0(fresh_wire_1141),
.PORT_ID_IN1(fresh_wire_1142),
.PORT_ID_OUT(fresh_wire_1143));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000020)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__233__DOLLAR__500$extendA(.PORT_ID_IN(fresh_wire_1144),
.PORT_ID_OUT(fresh_wire_1145));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000020)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__233__DOLLAR__500$op0(.PORT_ID_IN0(fresh_wire_1146),
.PORT_ID_IN1(fresh_wire_1147),
.PORT_ID_OUT(fresh_wire_1148));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000020)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__235__DOLLAR__501$extendA(.PORT_ID_IN(fresh_wire_1149),
.PORT_ID_OUT(fresh_wire_1150));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000020)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__235__DOLLAR__501$op0(.PORT_ID_IN0(fresh_wire_1151),
.PORT_ID_IN1(fresh_wire_1152),
.PORT_ID_OUT(fresh_wire_1153));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000020)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__242__DOLLAR__504$extendA(.PORT_ID_IN(fresh_wire_1154),
.PORT_ID_OUT(fresh_wire_1155));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000020)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__242__DOLLAR__504$op0(.PORT_ID_IN0(fresh_wire_1156),
.PORT_ID_IN1(fresh_wire_1157),
.PORT_ID_OUT(fresh_wire_1158));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__271__DOLLAR__521$op0(.PORT_ID_IN0(fresh_wire_1159),
.PORT_ID_IN1(fresh_wire_1160),
.PORT_ID_OUT(fresh_wire_1161));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__273__DOLLAR__525$op0(.PORT_ID_IN0(fresh_wire_1162),
.PORT_ID_IN1(fresh_wire_1163),
.PORT_ID_OUT(fresh_wire_1164));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__276__DOLLAR__534$op0(.PORT_ID_IN0(fresh_wire_1165),
.PORT_ID_IN1(fresh_wire_1166),
.PORT_ID_OUT(fresh_wire_1167));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__555$op0(.PORT_ID_IN0(fresh_wire_1168),
.PORT_ID_IN1(fresh_wire_1169),
.PORT_ID_OUT(fresh_wire_1170));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__207__DOLLAR__491$op0(.PORT_ID_IN0(fresh_wire_1171),
.PORT_ID_IN1(fresh_wire_1172),
.PORT_ID_OUT(fresh_wire_1173));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__466$op0(.PORT_ID_IN0(fresh_wire_1174),
.PORT_ID_IN1(fresh_wire_1175),
.PORT_ID_OUT(fresh_wire_1176));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__467$op0(.PORT_ID_IN0(fresh_wire_1177),
.PORT_ID_IN1(fresh_wire_1178),
.PORT_ID_OUT(fresh_wire_1179));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__469$op0(.PORT_ID_IN0(fresh_wire_1180),
.PORT_ID_IN1(fresh_wire_1181),
.PORT_ID_OUT(fresh_wire_1182));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__472$op0(.PORT_ID_IN0(fresh_wire_1183),
.PORT_ID_IN1(fresh_wire_1184),
.PORT_ID_OUT(fresh_wire_1185));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__176__DOLLAR__474$op0(.PORT_ID_IN0(fresh_wire_1186),
.PORT_ID_IN1(fresh_wire_1187),
.PORT_ID_OUT(fresh_wire_1188));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__192__DOLLAR__482$op0(.PORT_ID_IN0(fresh_wire_1189),
.PORT_ID_IN1(fresh_wire_1190),
.PORT_ID_OUT(fresh_wire_1191));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__193__DOLLAR__483$op0(.PORT_ID_IN0(fresh_wire_1192),
.PORT_ID_IN1(fresh_wire_1193),
.PORT_ID_OUT(fresh_wire_1194));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__196__DOLLAR__484$op0(.PORT_ID_IN0(fresh_wire_1195),
.PORT_ID_IN1(fresh_wire_1196),
.PORT_ID_OUT(fresh_wire_1197));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__207__DOLLAR__490$op0(.PORT_ID_IN0(fresh_wire_1198),
.PORT_ID_IN1(fresh_wire_1199),
.PORT_ID_OUT(fresh_wire_1200));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__228__DOLLAR__497$op0(.PORT_ID_IN0(fresh_wire_1201),
.PORT_ID_IN1(fresh_wire_1202),
.PORT_ID_OUT(fresh_wire_1203));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__229__DOLLAR__498$op0(.PORT_ID_IN0(fresh_wire_1204),
.PORT_ID_IN1(fresh_wire_1205),
.PORT_ID_OUT(fresh_wire_1206));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__268__DOLLAR__513$op0(.PORT_ID_IN0(fresh_wire_1207),
.PORT_ID_IN1(fresh_wire_1208),
.PORT_ID_OUT(fresh_wire_1209));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__268__DOLLAR__516$op0(.PORT_ID_IN0(fresh_wire_1210),
.PORT_ID_IN1(fresh_wire_1211),
.PORT_ID_OUT(fresh_wire_1212));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__273__DOLLAR__524$op0(.PORT_ID_IN0(fresh_wire_1213),
.PORT_ID_IN1(fresh_wire_1214),
.PORT_ID_OUT(fresh_wire_1215));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__285__DOLLAR__541$op0(.PORT_ID_IN0(fresh_wire_1216),
.PORT_ID_IN1(fresh_wire_1217),
.PORT_ID_OUT(fresh_wire_1218));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__309__DOLLAR__549$op0(.PORT_ID_IN0(fresh_wire_1219),
.PORT_ID_IN1(fresh_wire_1220),
.PORT_ID_OUT(fresh_wire_1221));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__556$op0(.PORT_ID_IN0(fresh_wire_1222),
.PORT_ID_IN1(fresh_wire_1223),
.PORT_ID_OUT(fresh_wire_1224));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__316__DOLLAR__558$op0(.PORT_ID_IN0(fresh_wire_1225),
.PORT_ID_IN1(fresh_wire_1226),
.PORT_ID_OUT(fresh_wire_1227));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__355__DOLLAR__568$op0(.PORT_ID_IN0(fresh_wire_1228),
.PORT_ID_IN1(fresh_wire_1229),
.PORT_ID_OUT(fresh_wire_1230));

	CELL_TYPE_UGE #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__ge__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__230__DOLLAR__499$op0(.PORT_ID_IN0(fresh_wire_1231),
.PORT_ID_IN1(fresh_wire_1232),
.PORT_ID_OUT(fresh_wire_1233));

	CELL_TYPE_UGE #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__ge__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__239__DOLLAR__503$op0(.PORT_ID_IN0(fresh_wire_1234),
.PORT_ID_IN1(fresh_wire_1235),
.PORT_ID_OUT(fresh_wire_1236));

	CELL_TYPE_UGE #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__ge__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__276__DOLLAR__535$op0(.PORT_ID_IN0(fresh_wire_1237),
.PORT_ID_IN1(fresh_wire_1238),
.PORT_ID_OUT(fresh_wire_1239));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__468$aRed(.PORT_ID_IN(fresh_wire_1240),
.PORT_ID_OUT(fresh_wire_1241));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__468$andOps(.PORT_ID_IN0(fresh_wire_1242),
.PORT_ID_IN1(fresh_wire_1243),
.PORT_ID_OUT(fresh_wire_1244));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__468$bRed(.PORT_ID_IN(fresh_wire_1245),
.PORT_ID_OUT(fresh_wire_1246));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__470$aRed(.PORT_ID_IN(fresh_wire_1247),
.PORT_ID_OUT(fresh_wire_1248));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__470$andOps(.PORT_ID_IN0(fresh_wire_1249),
.PORT_ID_IN1(fresh_wire_1250),
.PORT_ID_OUT(fresh_wire_1251));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__470$bRed(.PORT_ID_IN(fresh_wire_1252),
.PORT_ID_OUT(fresh_wire_1253));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__473$aRed(.PORT_ID_IN(fresh_wire_1254),
.PORT_ID_OUT(fresh_wire_1255));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__473$andOps(.PORT_ID_IN0(fresh_wire_1256),
.PORT_ID_IN1(fresh_wire_1257),
.PORT_ID_OUT(fresh_wire_1258));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__175__DOLLAR__473$bRed(.PORT_ID_IN(fresh_wire_1259),
.PORT_ID_OUT(fresh_wire_1260));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__268__DOLLAR__515$aRed(.PORT_ID_IN(fresh_wire_1261),
.PORT_ID_OUT(fresh_wire_1262));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__268__DOLLAR__515$andOps(.PORT_ID_IN0(fresh_wire_1263),
.PORT_ID_IN1(fresh_wire_1264),
.PORT_ID_OUT(fresh_wire_1265));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__268__DOLLAR__517$aRed(.PORT_ID_IN(fresh_wire_1266),
.PORT_ID_OUT(fresh_wire_1267));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__268__DOLLAR__517$andOps(.PORT_ID_IN0(fresh_wire_1268),
.PORT_ID_IN1(fresh_wire_1269),
.PORT_ID_OUT(fresh_wire_1270));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__268__DOLLAR__517$bRed(.PORT_ID_IN(fresh_wire_1271),
.PORT_ID_OUT(fresh_wire_1272));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__271__DOLLAR__520$aRed(.PORT_ID_IN(fresh_wire_1273),
.PORT_ID_OUT(fresh_wire_1274));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__271__DOLLAR__520$andOps(.PORT_ID_IN0(fresh_wire_1275),
.PORT_ID_IN1(fresh_wire_1276),
.PORT_ID_OUT(fresh_wire_1277));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__271__DOLLAR__523$aRed(.PORT_ID_IN(fresh_wire_1278),
.PORT_ID_OUT(fresh_wire_1279));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__271__DOLLAR__523$andOps(.PORT_ID_IN0(fresh_wire_1280),
.PORT_ID_IN1(fresh_wire_1281),
.PORT_ID_OUT(fresh_wire_1282));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__271__DOLLAR__523$bRed(.PORT_ID_IN(fresh_wire_1283),
.PORT_ID_OUT(fresh_wire_1284));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__276__DOLLAR__536$aRed(.PORT_ID_IN(fresh_wire_1285),
.PORT_ID_OUT(fresh_wire_1286));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__276__DOLLAR__536$andOps(.PORT_ID_IN0(fresh_wire_1287),
.PORT_ID_IN1(fresh_wire_1288),
.PORT_ID_OUT(fresh_wire_1289));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__276__DOLLAR__536$bRed(.PORT_ID_IN(fresh_wire_1290),
.PORT_ID_OUT(fresh_wire_1291));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__277__DOLLAR__539$andOps(.PORT_ID_IN0(fresh_wire_1292),
.PORT_ID_IN1(fresh_wire_1293),
.PORT_ID_OUT(fresh_wire_1294));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__277__DOLLAR__539$bRed(.PORT_ID_IN(fresh_wire_1295),
.PORT_ID_OUT(fresh_wire_1296));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__285__DOLLAR__543$aRed(.PORT_ID_IN(fresh_wire_1297),
.PORT_ID_OUT(fresh_wire_1298));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__285__DOLLAR__543$andOps(.PORT_ID_IN0(fresh_wire_1299),
.PORT_ID_IN1(fresh_wire_1300),
.PORT_ID_OUT(fresh_wire_1301));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__552$aRed(.PORT_ID_IN(fresh_wire_1302),
.PORT_ID_OUT(fresh_wire_1303));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__552$andOps(.PORT_ID_IN0(fresh_wire_1304),
.PORT_ID_IN1(fresh_wire_1305),
.PORT_ID_OUT(fresh_wire_1306));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__552$bRed(.PORT_ID_IN(fresh_wire_1307),
.PORT_ID_OUT(fresh_wire_1308));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__554$aRed(.PORT_ID_IN(fresh_wire_1309),
.PORT_ID_OUT(fresh_wire_1310));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__554$andOps(.PORT_ID_IN0(fresh_wire_1311),
.PORT_ID_IN1(fresh_wire_1312),
.PORT_ID_OUT(fresh_wire_1313));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__554$bRed(.PORT_ID_IN(fresh_wire_1314),
.PORT_ID_OUT(fresh_wire_1315));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__557$aRed(.PORT_ID_IN(fresh_wire_1316),
.PORT_ID_OUT(fresh_wire_1317));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__557$andOps(.PORT_ID_IN0(fresh_wire_1318),
.PORT_ID_IN1(fresh_wire_1319),
.PORT_ID_OUT(fresh_wire_1320));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__312__DOLLAR__557$bRed(.PORT_ID_IN(fresh_wire_1321),
.PORT_ID_OUT(fresh_wire_1322));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__316__DOLLAR__560$aRed(.PORT_ID_IN(fresh_wire_1323),
.PORT_ID_OUT(fresh_wire_1324));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__316__DOLLAR__560$andOps(.PORT_ID_IN0(fresh_wire_1325),
.PORT_ID_IN1(fresh_wire_1326),
.PORT_ID_OUT(fresh_wire_1327));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_or__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__344__DOLLAR__565$bRed(.PORT_ID_IN(fresh_wire_1328),
.PORT_ID_OUT(fresh_wire_1329));

	CELL_TYPE_OR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__logic_or__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__344__DOLLAR__565$orOps(.PORT_ID_IN0(fresh_wire_1330),
.PORT_ID_IN1(fresh_wire_1331),
.PORT_ID_OUT(fresh_wire_1332));

	CELL_TYPE_ULT #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__lt__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__250__DOLLAR__507$op0(.PORT_ID_IN0(fresh_wire_1333),
.PORT_ID_IN1(fresh_wire_1334),
.PORT_ID_OUT(fresh_wire_1335));

	CELL_TYPE_ULT #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__lt__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__271__DOLLAR__522$op0(.PORT_ID_IN0(fresh_wire_1336),
.PORT_ID_IN1(fresh_wire_1337),
.PORT_ID_OUT(fresh_wire_1338));

	CELL_TYPE_NOT #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__not__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__171__DOLLAR__465$op0(.PORT_ID_IN(fresh_wire_1339),
.PORT_ID_OUT(fresh_wire_1340));

	CELL_TYPE_REG #(.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3712$reg0(.PORT_ID_CLK(fresh_wire_1343),
.PORT_ID_IN(fresh_wire_1341),
.PORT_ID_OUT(fresh_wire_1342));

	CELL_TYPE_REG #(.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(2'hx),
.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3713$reg0(.PORT_ID_CLK(fresh_wire_1346),
.PORT_ID_IN(fresh_wire_1344),
.PORT_ID_OUT(fresh_wire_1345));

	CELL_TYPE_REG #(.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(2'hx),
.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3714$reg0(.PORT_ID_CLK(fresh_wire_1349),
.PORT_ID_IN(fresh_wire_1347),
.PORT_ID_OUT(fresh_wire_1348));

	CELL_TYPE_REG #(.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(16'hxxxx),
.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3716$reg0(.PORT_ID_CLK(fresh_wire_1352),
.PORT_ID_IN(fresh_wire_1350),
.PORT_ID_OUT(fresh_wire_1351));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3718$reg0(.PORT_ID_ARST(fresh_wire_1356),
.PORT_ID_CLK(fresh_wire_1355),
.PORT_ID_IN(fresh_wire_1353),
.PORT_ID_OUT(fresh_wire_1354));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3719$reg0(.PORT_ID_ARST(fresh_wire_1360),
.PORT_ID_CLK(fresh_wire_1359),
.PORT_ID_IN(fresh_wire_1357),
.PORT_ID_OUT(fresh_wire_1358));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3720$reg0(.PORT_ID_ARST(fresh_wire_1364),
.PORT_ID_CLK(fresh_wire_1363),
.PORT_ID_IN(fresh_wire_1361),
.PORT_ID_OUT(fresh_wire_1362));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3721$reg0(.PORT_ID_ARST(fresh_wire_1368),
.PORT_ID_CLK(fresh_wire_1367),
.PORT_ID_IN(fresh_wire_1365),
.PORT_ID_OUT(fresh_wire_1366));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3722$reg0(.PORT_ID_ARST(fresh_wire_1372),
.PORT_ID_CLK(fresh_wire_1371),
.PORT_ID_IN(fresh_wire_1369),
.PORT_ID_OUT(fresh_wire_1370));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(2'h0),
.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3723$reg0(.PORT_ID_ARST(fresh_wire_1376),
.PORT_ID_CLK(fresh_wire_1375),
.PORT_ID_IN(fresh_wire_1373),
.PORT_ID_OUT(fresh_wire_1374));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(16'h0000),
.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3724$reg0(.PORT_ID_ARST(fresh_wire_1380),
.PORT_ID_CLK(fresh_wire_1379),
.PORT_ID_IN(fresh_wire_1377),
.PORT_ID_OUT(fresh_wire_1378));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(16'h0000),
.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3725$reg0(.PORT_ID_ARST(fresh_wire_1384),
.PORT_ID_CLK(fresh_wire_1383),
.PORT_ID_IN(fresh_wire_1381),
.PORT_ID_OUT(fresh_wire_1382));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(16'h0000),
.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3726$reg0(.PORT_ID_ARST(fresh_wire_1388),
.PORT_ID_CLK(fresh_wire_1387),
.PORT_ID_IN(fresh_wire_1385),
.PORT_ID_OUT(fresh_wire_1386));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(16'h0000),
.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3727$reg0(.PORT_ID_ARST(fresh_wire_1392),
.PORT_ID_CLK(fresh_wire_1391),
.PORT_ID_IN(fresh_wire_1389),
.PORT_ID_OUT(fresh_wire_1390));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3728$reg0(.PORT_ID_ARST(fresh_wire_1396),
.PORT_ID_CLK(fresh_wire_1395),
.PORT_ID_IN(fresh_wire_1393),
.PORT_ID_OUT(fresh_wire_1394));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3729$reg0(.PORT_ID_ARST(fresh_wire_1400),
.PORT_ID_CLK(fresh_wire_1399),
.PORT_ID_IN(fresh_wire_1397),
.PORT_ID_OUT(fresh_wire_1398));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procdff__DOLLAR__3730$reg0(.PORT_ID_ARST(fresh_wire_1404),
.PORT_ID_CLK(fresh_wire_1403),
.PORT_ID_IN(fresh_wire_1401),
.PORT_ID_OUT(fresh_wire_1402));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2788$mux0(.PORT_ID_IN0(fresh_wire_1405),
.PORT_ID_IN1(fresh_wire_1406),
.PORT_ID_OUT(fresh_wire_1407),
.PORT_ID_SEL(fresh_wire_1408));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2865$mux0(.PORT_ID_IN0(fresh_wire_1409),
.PORT_ID_IN1(fresh_wire_1410),
.PORT_ID_OUT(fresh_wire_1411),
.PORT_ID_SEL(fresh_wire_1412));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2867$mux0(.PORT_ID_IN0(fresh_wire_1413),
.PORT_ID_IN1(fresh_wire_1414),
.PORT_ID_OUT(fresh_wire_1415),
.PORT_ID_SEL(fresh_wire_1416));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2877$mux0(.PORT_ID_IN0(fresh_wire_1417),
.PORT_ID_IN1(fresh_wire_1418),
.PORT_ID_OUT(fresh_wire_1419),
.PORT_ID_SEL(fresh_wire_1420));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2879$mux0(.PORT_ID_IN0(fresh_wire_1421),
.PORT_ID_IN1(fresh_wire_1422),
.PORT_ID_OUT(fresh_wire_1423),
.PORT_ID_SEL(fresh_wire_1424));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2888$mux0(.PORT_ID_IN0(fresh_wire_1425),
.PORT_ID_IN1(fresh_wire_1426),
.PORT_ID_OUT(fresh_wire_1427),
.PORT_ID_SEL(fresh_wire_1428));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2898$mux0(.PORT_ID_IN0(fresh_wire_1429),
.PORT_ID_IN1(fresh_wire_1430),
.PORT_ID_OUT(fresh_wire_1431),
.PORT_ID_SEL(fresh_wire_1432));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2904$mux0(.PORT_ID_IN0(fresh_wire_1433),
.PORT_ID_IN1(fresh_wire_1434),
.PORT_ID_OUT(fresh_wire_1435),
.PORT_ID_SEL(fresh_wire_1436));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2907$mux0(.PORT_ID_IN0(fresh_wire_1437),
.PORT_ID_IN1(fresh_wire_1438),
.PORT_ID_OUT(fresh_wire_1439),
.PORT_ID_SEL(fresh_wire_1440));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2909$mux0(.PORT_ID_IN0(fresh_wire_1441),
.PORT_ID_IN1(fresh_wire_1442),
.PORT_ID_OUT(fresh_wire_1443),
.PORT_ID_SEL(fresh_wire_1444));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2919$mux0(.PORT_ID_IN0(fresh_wire_1445),
.PORT_ID_IN1(fresh_wire_1446),
.PORT_ID_OUT(fresh_wire_1447),
.PORT_ID_SEL(fresh_wire_1448));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2923$mux0(.PORT_ID_IN0(fresh_wire_1449),
.PORT_ID_IN1(fresh_wire_1450),
.PORT_ID_OUT(fresh_wire_1451),
.PORT_ID_SEL(fresh_wire_1452));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2925$mux0(.PORT_ID_IN0(fresh_wire_1453),
.PORT_ID_IN1(fresh_wire_1454),
.PORT_ID_OUT(fresh_wire_1455),
.PORT_ID_SEL(fresh_wire_1456));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2931$mux0(.PORT_ID_IN0(fresh_wire_1457),
.PORT_ID_IN1(fresh_wire_1458),
.PORT_ID_OUT(fresh_wire_1459),
.PORT_ID_SEL(fresh_wire_1460));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2934$mux0(.PORT_ID_IN0(fresh_wire_1461),
.PORT_ID_IN1(fresh_wire_1462),
.PORT_ID_OUT(fresh_wire_1463),
.PORT_ID_SEL(fresh_wire_1464));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2936$mux0(.PORT_ID_IN0(fresh_wire_1465),
.PORT_ID_IN1(fresh_wire_1466),
.PORT_ID_OUT(fresh_wire_1467),
.PORT_ID_SEL(fresh_wire_1468));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2946$mux0(.PORT_ID_IN0(fresh_wire_1469),
.PORT_ID_IN1(fresh_wire_1470),
.PORT_ID_OUT(fresh_wire_1471),
.PORT_ID_SEL(fresh_wire_1472));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2952$mux0(.PORT_ID_IN0(fresh_wire_1473),
.PORT_ID_IN1(fresh_wire_1474),
.PORT_ID_OUT(fresh_wire_1475),
.PORT_ID_SEL(fresh_wire_1476));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2955$mux0(.PORT_ID_IN0(fresh_wire_1477),
.PORT_ID_IN1(fresh_wire_1478),
.PORT_ID_OUT(fresh_wire_1479),
.PORT_ID_SEL(fresh_wire_1480));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2957$mux0(.PORT_ID_IN0(fresh_wire_1481),
.PORT_ID_IN1(fresh_wire_1482),
.PORT_ID_OUT(fresh_wire_1483),
.PORT_ID_SEL(fresh_wire_1484));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2967$mux0(.PORT_ID_IN0(fresh_wire_1485),
.PORT_ID_IN1(fresh_wire_1486),
.PORT_ID_OUT(fresh_wire_1487),
.PORT_ID_SEL(fresh_wire_1488));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2971$mux0(.PORT_ID_IN0(fresh_wire_1489),
.PORT_ID_IN1(fresh_wire_1490),
.PORT_ID_OUT(fresh_wire_1491),
.PORT_ID_SEL(fresh_wire_1492));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2973$mux0(.PORT_ID_IN0(fresh_wire_1493),
.PORT_ID_IN1(fresh_wire_1494),
.PORT_ID_OUT(fresh_wire_1495),
.PORT_ID_SEL(fresh_wire_1496));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2979$mux0(.PORT_ID_IN0(fresh_wire_1497),
.PORT_ID_IN1(fresh_wire_1498),
.PORT_ID_OUT(fresh_wire_1499),
.PORT_ID_SEL(fresh_wire_1500));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2982$mux0(.PORT_ID_IN0(fresh_wire_1501),
.PORT_ID_IN1(fresh_wire_1502),
.PORT_ID_OUT(fresh_wire_1503),
.PORT_ID_SEL(fresh_wire_1504));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2984$mux0(.PORT_ID_IN0(fresh_wire_1505),
.PORT_ID_IN1(fresh_wire_1506),
.PORT_ID_OUT(fresh_wire_1507),
.PORT_ID_SEL(fresh_wire_1508));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2993$mux0(.PORT_ID_IN0(fresh_wire_1509),
.PORT_ID_IN1(fresh_wire_1510),
.PORT_ID_OUT(fresh_wire_1511),
.PORT_ID_SEL(fresh_wire_1512));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2997$mux0(.PORT_ID_IN0(fresh_wire_1513),
.PORT_ID_IN1(fresh_wire_1514),
.PORT_ID_OUT(fresh_wire_1515),
.PORT_ID_SEL(fresh_wire_1516));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__2999$mux0(.PORT_ID_IN0(fresh_wire_1517),
.PORT_ID_IN1(fresh_wire_1518),
.PORT_ID_OUT(fresh_wire_1519),
.PORT_ID_SEL(fresh_wire_1520));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3013$mux0(.PORT_ID_IN0(fresh_wire_1521),
.PORT_ID_IN1(fresh_wire_1522),
.PORT_ID_OUT(fresh_wire_1523),
.PORT_ID_SEL(fresh_wire_1524));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3015$mux0(.PORT_ID_IN0(fresh_wire_1525),
.PORT_ID_IN1(fresh_wire_1526),
.PORT_ID_OUT(fresh_wire_1527),
.PORT_ID_SEL(fresh_wire_1528));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3017$mux0(.PORT_ID_IN0(fresh_wire_1529),
.PORT_ID_IN1(fresh_wire_1530),
.PORT_ID_OUT(fresh_wire_1531),
.PORT_ID_SEL(fresh_wire_1532));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3033$mux0(.PORT_ID_IN0(fresh_wire_1533),
.PORT_ID_IN1(fresh_wire_1534),
.PORT_ID_OUT(fresh_wire_1535),
.PORT_ID_SEL(fresh_wire_1536));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3035$mux0(.PORT_ID_IN0(fresh_wire_1537),
.PORT_ID_IN1(fresh_wire_1538),
.PORT_ID_OUT(fresh_wire_1539),
.PORT_ID_SEL(fresh_wire_1540));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3038$mux0(.PORT_ID_IN0(fresh_wire_1541),
.PORT_ID_IN1(fresh_wire_1542),
.PORT_ID_OUT(fresh_wire_1543),
.PORT_ID_SEL(fresh_wire_1544));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3057$mux0(.PORT_ID_IN0(fresh_wire_1545),
.PORT_ID_IN1(fresh_wire_1546),
.PORT_ID_OUT(fresh_wire_1547),
.PORT_ID_SEL(fresh_wire_1548));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3059$mux0(.PORT_ID_IN0(fresh_wire_1549),
.PORT_ID_IN1(fresh_wire_1550),
.PORT_ID_OUT(fresh_wire_1551),
.PORT_ID_SEL(fresh_wire_1552));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3069$mux0(.PORT_ID_IN0(fresh_wire_1553),
.PORT_ID_IN1(fresh_wire_1554),
.PORT_ID_OUT(fresh_wire_1555),
.PORT_ID_SEL(fresh_wire_1556));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3072$mux0(.PORT_ID_IN0(fresh_wire_1557),
.PORT_ID_IN1(fresh_wire_1558),
.PORT_ID_OUT(fresh_wire_1559),
.PORT_ID_SEL(fresh_wire_1560));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__procmux__DOLLAR__3074$mux0(.PORT_ID_IN0(fresh_wire_1561),
.PORT_ID_IN1(fresh_wire_1562),
.PORT_ID_OUT(fresh_wire_1563),
.PORT_ID_SEL(fresh_wire_1564));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000020)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__sub__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__244__DOLLAR__505$extendA(.PORT_ID_IN(fresh_wire_1565),
.PORT_ID_OUT(fresh_wire_1566));

	CELL_TYPE_SUB #(.PARAM_WIDTH(32'h00000020)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__sub__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__244__DOLLAR__505$op0(.PORT_ID_IN0(fresh_wire_1567),
.PORT_ID_IN1(fresh_wire_1568),
.PORT_ID_OUT(fresh_wire_1569));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000020)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__ternary__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__176__DOLLAR__475$mux0(.PORT_ID_IN0(fresh_wire_1570),
.PORT_ID_IN1(fresh_wire_1571),
.PORT_ID_OUT(fresh_wire_1572),
.PORT_ID_SEL(fresh_wire_1573));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__ternary__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__273__DOLLAR__526$mux0(.PORT_ID_IN0(fresh_wire_1574),
.PORT_ID_IN1(fresh_wire_1575),
.PORT_ID_OUT(fresh_wire_1576),
.PORT_ID_SEL(fresh_wire_1577));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__ternary__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__273__DOLLAR__526__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(.PORT_ID_OUT(fresh_wire_1578));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$__DOLLAR__ternary__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__linebuffer_control_unq1__DOT__v__COLON__355__DOLLAR__569$mux0(.PORT_ID_IN0(fresh_wire_1579),
.PORT_ID_IN1(fresh_wire_1580),
.PORT_ID_OUT(fresh_wire_1581),
.PORT_ID_SEL(fresh_wire_1582));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__101__DOLLAR__314$op0(.PORT_ID_IN0(fresh_wire_1583),
.PORT_ID_IN1(fresh_wire_1584),
.PORT_ID_OUT(fresh_wire_1585));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__100__DOLLAR__310$op0(.PORT_ID_IN0(fresh_wire_1586),
.PORT_ID_IN1(fresh_wire_1587),
.PORT_ID_OUT(fresh_wire_1588));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__100__DOLLAR__311$op0(.PORT_ID_IN0(fresh_wire_1589),
.PORT_ID_IN1(fresh_wire_1590),
.PORT_ID_OUT(fresh_wire_1591));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__103__DOLLAR__316$op0(.PORT_ID_IN0(fresh_wire_1592),
.PORT_ID_IN1(fresh_wire_1593),
.PORT_ID_OUT(fresh_wire_1594));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__128__DOLLAR__345$op0(.PORT_ID_IN0(fresh_wire_1595),
.PORT_ID_IN1(fresh_wire_1596),
.PORT_ID_OUT(fresh_wire_1597));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__150__DOLLAR__379$op0(.PORT_ID_IN0(fresh_wire_1598),
.PORT_ID_IN1(fresh_wire_1599),
.PORT_ID_OUT(fresh_wire_1600));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__157__DOLLAR__381$op0(.PORT_ID_IN0(fresh_wire_1601),
.PORT_ID_IN1(fresh_wire_1602),
.PORT_ID_OUT(fresh_wire_1603));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__158__DOLLAR__382$op0(.PORT_ID_IN0(fresh_wire_1604),
.PORT_ID_IN1(fresh_wire_1605),
.PORT_ID_OUT(fresh_wire_1606));

	CELL_TYPE_UGE #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__ge__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__126__DOLLAR__341$op0(.PORT_ID_IN0(fresh_wire_1607),
.PORT_ID_IN1(fresh_wire_1608),
.PORT_ID_OUT(fresh_wire_1609));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__100__DOLLAR__312$aRed(.PORT_ID_IN(fresh_wire_1610),
.PORT_ID_OUT(fresh_wire_1611));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__100__DOLLAR__312$andOps(.PORT_ID_IN0(fresh_wire_1612),
.PORT_ID_IN1(fresh_wire_1613),
.PORT_ID_OUT(fresh_wire_1614));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__100__DOLLAR__312$bRed(.PORT_ID_IN(fresh_wire_1615),
.PORT_ID_OUT(fresh_wire_1616));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__100__DOLLAR__313$andOps(.PORT_ID_IN0(fresh_wire_1617),
.PORT_ID_IN1(fresh_wire_1618),
.PORT_ID_OUT(fresh_wire_1619));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__100__DOLLAR__313$bRed(.PORT_ID_IN(fresh_wire_1620),
.PORT_ID_OUT(fresh_wire_1621));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__103__DOLLAR__317$andOps(.PORT_ID_IN0(fresh_wire_1622),
.PORT_ID_IN1(fresh_wire_1623),
.PORT_ID_OUT(fresh_wire_1624));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__103__DOLLAR__317$bRed(.PORT_ID_IN(fresh_wire_1625),
.PORT_ID_OUT(fresh_wire_1626));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__125__DOLLAR__340$andOps(.PORT_ID_IN0(fresh_wire_1627),
.PORT_ID_IN1(fresh_wire_1628),
.PORT_ID_OUT(fresh_wire_1629));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__125__DOLLAR__340$bRed(.PORT_ID_IN(fresh_wire_1630),
.PORT_ID_OUT(fresh_wire_1631));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__127__DOLLAR__344$andOps(.PORT_ID_IN0(fresh_wire_1632),
.PORT_ID_IN1(fresh_wire_1633),
.PORT_ID_OUT(fresh_wire_1634));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__127__DOLLAR__344$bRed(.PORT_ID_IN(fresh_wire_1635),
.PORT_ID_OUT(fresh_wire_1636));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(2'h0),
.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__procdff__DOLLAR__3739$reg0(.PORT_ID_ARST(fresh_wire_1640),
.PORT_ID_CLK(fresh_wire_1639),
.PORT_ID_IN(fresh_wire_1637),
.PORT_ID_OUT(fresh_wire_1638));

	CELL_TYPE_REG #(.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(48'hxxxxxxxxxxxx),
.PARAM_WIDTH(32'h00000030)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__procdff__DOLLAR__3740$reg0(.PORT_ID_CLK(fresh_wire_1643),
.PORT_ID_IN(fresh_wire_1641),
.PORT_ID_OUT(fresh_wire_1642));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3178$mux0(.PORT_ID_IN0(fresh_wire_1644),
.PORT_ID_IN1(fresh_wire_1645),
.PORT_ID_OUT(fresh_wire_1646),
.PORT_ID_SEL(fresh_wire_1647));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3181$mux0(.PORT_ID_IN0(fresh_wire_1648),
.PORT_ID_IN1(fresh_wire_1649),
.PORT_ID_OUT(fresh_wire_1650),
.PORT_ID_SEL(fresh_wire_1651));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3199$mux0(.PORT_ID_IN0(fresh_wire_1652),
.PORT_ID_IN1(fresh_wire_1653),
.PORT_ID_OUT(fresh_wire_1654),
.PORT_ID_SEL(fresh_wire_1655));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3202$mux0(.PORT_ID_IN0(fresh_wire_1656),
.PORT_ID_IN1(fresh_wire_1657),
.PORT_ID_OUT(fresh_wire_1658),
.PORT_ID_SEL(fresh_wire_1659));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000020)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3211$mux0(.PORT_ID_IN0(fresh_wire_1660),
.PORT_ID_IN1(fresh_wire_1661),
.PORT_ID_OUT(fresh_wire_1662),
.PORT_ID_SEL(fresh_wire_1663));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000020)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3214$mux0(.PORT_ID_IN0(fresh_wire_1664),
.PORT_ID_IN1(fresh_wire_1665),
.PORT_ID_OUT(fresh_wire_1666),
.PORT_ID_SEL(fresh_wire_1667));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000020)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3217$mux0(.PORT_ID_IN0(fresh_wire_1668),
.PORT_ID_IN1(fresh_wire_1669),
.PORT_ID_OUT(fresh_wire_1670),
.PORT_ID_SEL(fresh_wire_1671));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000020)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3219$mux0(.PORT_ID_IN0(fresh_wire_1672),
.PORT_ID_IN1(fresh_wire_1673),
.PORT_ID_OUT(fresh_wire_1674),
.PORT_ID_SEL(fresh_wire_1675));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000020)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3223$mux0(.PORT_ID_IN0(fresh_wire_1676),
.PORT_ID_IN1(fresh_wire_1677),
.PORT_ID_OUT(fresh_wire_1678),
.PORT_ID_SEL(fresh_wire_1679));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000020)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3226$mux0(.PORT_ID_IN0(fresh_wire_1680),
.PORT_ID_IN1(fresh_wire_1681),
.PORT_ID_OUT(fresh_wire_1682),
.PORT_ID_SEL(fresh_wire_1683));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000020)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__procmux__DOLLAR__3228$mux0(.PORT_ID_IN0(fresh_wire_1684),
.PORT_ID_IN1(fresh_wire_1685),
.PORT_ID_OUT(fresh_wire_1686),
.PORT_ID_SEL(fresh_wire_1687));

	CELL_TYPE_SUB #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__sub__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__104__DOLLAR__318$op0(.PORT_ID_IN0(fresh_wire_1688),
.PORT_ID_IN1(fresh_wire_1689),
.PORT_ID_OUT(fresh_wire_1690));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$input_sr$__DOLLAR__sub__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__input_sr_unq1__DOT__v__COLON__110__DOLLAR__326__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(.PORT_ID_OUT(fresh_wire_1691));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__103__DOLLAR__747$op0(.PORT_ID_IN0(fresh_wire_1692),
.PORT_ID_IN1(fresh_wire_1693),
.PORT_ID_OUT(fresh_wire_1694));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__106__DOLLAR__751$op0(.PORT_ID_IN0(fresh_wire_1695),
.PORT_ID_IN1(fresh_wire_1696),
.PORT_ID_OUT(fresh_wire_1697));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__102__DOLLAR__744$op0(.PORT_ID_IN0(fresh_wire_1698),
.PORT_ID_IN1(fresh_wire_1699),
.PORT_ID_OUT(fresh_wire_1700));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__102__DOLLAR__745$op0(.PORT_ID_IN0(fresh_wire_1701),
.PORT_ID_IN1(fresh_wire_1702),
.PORT_ID_OUT(fresh_wire_1703));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__105__DOLLAR__748$op0(.PORT_ID_IN0(fresh_wire_1704),
.PORT_ID_IN1(fresh_wire_1705),
.PORT_ID_OUT(fresh_wire_1706));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__108__DOLLAR__753$op0(.PORT_ID_IN0(fresh_wire_1707),
.PORT_ID_IN1(fresh_wire_1708),
.PORT_ID_OUT(fresh_wire_1709));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__120__DOLLAR__760$op0(.PORT_ID_IN0(fresh_wire_1710),
.PORT_ID_IN1(fresh_wire_1711),
.PORT_ID_OUT(fresh_wire_1712));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__120__DOLLAR__761$op0(.PORT_ID_IN0(fresh_wire_1713),
.PORT_ID_IN1(fresh_wire_1714),
.PORT_ID_OUT(fresh_wire_1715));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__133__DOLLAR__784$op0(.PORT_ID_IN0(fresh_wire_1716),
.PORT_ID_IN1(fresh_wire_1717),
.PORT_ID_OUT(fresh_wire_1718));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__135__DOLLAR__785$op0(.PORT_ID_IN0(fresh_wire_1719),
.PORT_ID_IN1(fresh_wire_1720),
.PORT_ID_OUT(fresh_wire_1721));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__137__DOLLAR__786$op0(.PORT_ID_IN0(fresh_wire_1722),
.PORT_ID_IN1(fresh_wire_1723),
.PORT_ID_OUT(fresh_wire_1724));

	CELL_TYPE_UGE #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__ge__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__121__DOLLAR__765$op0(.PORT_ID_IN0(fresh_wire_1725),
.PORT_ID_IN1(fresh_wire_1726),
.PORT_ID_OUT(fresh_wire_1727));

	CELL_TYPE_UGE #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__ge__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__123__DOLLAR__771$op0(.PORT_ID_IN0(fresh_wire_1728),
.PORT_ID_IN1(fresh_wire_1729),
.PORT_ID_OUT(fresh_wire_1730));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__102__DOLLAR__746$aRed(.PORT_ID_IN(fresh_wire_1731),
.PORT_ID_OUT(fresh_wire_1732));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__102__DOLLAR__746$andOps(.PORT_ID_IN0(fresh_wire_1733),
.PORT_ID_IN1(fresh_wire_1734),
.PORT_ID_OUT(fresh_wire_1735));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__102__DOLLAR__746$bRed(.PORT_ID_IN(fresh_wire_1736),
.PORT_ID_OUT(fresh_wire_1737));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__105__DOLLAR__750$aRed(.PORT_ID_IN(fresh_wire_1738),
.PORT_ID_OUT(fresh_wire_1739));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__105__DOLLAR__750$andOps(.PORT_ID_IN0(fresh_wire_1740),
.PORT_ID_IN1(fresh_wire_1741),
.PORT_ID_OUT(fresh_wire_1742));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__105__DOLLAR__750$bRed(.PORT_ID_IN(fresh_wire_1743),
.PORT_ID_OUT(fresh_wire_1744));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__108__DOLLAR__754$aRed(.PORT_ID_IN(fresh_wire_1745),
.PORT_ID_OUT(fresh_wire_1746));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__108__DOLLAR__754$andOps(.PORT_ID_IN0(fresh_wire_1747),
.PORT_ID_IN1(fresh_wire_1748),
.PORT_ID_OUT(fresh_wire_1749));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__108__DOLLAR__754$bRed(.PORT_ID_IN(fresh_wire_1750),
.PORT_ID_OUT(fresh_wire_1751));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__110__DOLLAR__757$aRed(.PORT_ID_IN(fresh_wire_1752),
.PORT_ID_OUT(fresh_wire_1753));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__110__DOLLAR__757$andOps(.PORT_ID_IN0(fresh_wire_1754),
.PORT_ID_IN1(fresh_wire_1755),
.PORT_ID_OUT(fresh_wire_1756));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__110__DOLLAR__757$bRed(.PORT_ID_IN(fresh_wire_1757),
.PORT_ID_OUT(fresh_wire_1758));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__120__DOLLAR__762$aRed(.PORT_ID_IN(fresh_wire_1759),
.PORT_ID_OUT(fresh_wire_1760));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__120__DOLLAR__762$andOps(.PORT_ID_IN0(fresh_wire_1761),
.PORT_ID_IN1(fresh_wire_1762),
.PORT_ID_OUT(fresh_wire_1763));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__120__DOLLAR__762$bRed(.PORT_ID_IN(fresh_wire_1764),
.PORT_ID_OUT(fresh_wire_1765));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__120__DOLLAR__764$aRed(.PORT_ID_IN(fresh_wire_1766),
.PORT_ID_OUT(fresh_wire_1767));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__120__DOLLAR__764$andOps(.PORT_ID_IN0(fresh_wire_1768),
.PORT_ID_IN1(fresh_wire_1769),
.PORT_ID_OUT(fresh_wire_1770));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__120__DOLLAR__764$bRed(.PORT_ID_IN(fresh_wire_1771),
.PORT_ID_OUT(fresh_wire_1772));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__122__DOLLAR__768$aRed(.PORT_ID_IN(fresh_wire_1773),
.PORT_ID_OUT(fresh_wire_1774));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__122__DOLLAR__768$andOps(.PORT_ID_IN0(fresh_wire_1775),
.PORT_ID_IN1(fresh_wire_1776),
.PORT_ID_OUT(fresh_wire_1777));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__122__DOLLAR__768$bRed(.PORT_ID_IN(fresh_wire_1778),
.PORT_ID_OUT(fresh_wire_1779));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__122__DOLLAR__770$aRed(.PORT_ID_IN(fresh_wire_1780),
.PORT_ID_OUT(fresh_wire_1781));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__122__DOLLAR__770$andOps(.PORT_ID_IN0(fresh_wire_1782),
.PORT_ID_IN1(fresh_wire_1783),
.PORT_ID_OUT(fresh_wire_1784));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__122__DOLLAR__770$bRed(.PORT_ID_IN(fresh_wire_1785),
.PORT_ID_OUT(fresh_wire_1786));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__124__DOLLAR__776$aRed(.PORT_ID_IN(fresh_wire_1787),
.PORT_ID_OUT(fresh_wire_1788));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__124__DOLLAR__776$andOps(.PORT_ID_IN0(fresh_wire_1789),
.PORT_ID_IN1(fresh_wire_1790),
.PORT_ID_OUT(fresh_wire_1791));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__124__DOLLAR__776$bRed(.PORT_ID_IN(fresh_wire_1792),
.PORT_ID_OUT(fresh_wire_1793));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__126__DOLLAR__781$aRed(.PORT_ID_IN(fresh_wire_1794),
.PORT_ID_OUT(fresh_wire_1795));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__126__DOLLAR__781$andOps(.PORT_ID_IN0(fresh_wire_1796),
.PORT_ID_IN1(fresh_wire_1797),
.PORT_ID_OUT(fresh_wire_1798));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__126__DOLLAR__781$bRed(.PORT_ID_IN(fresh_wire_1799),
.PORT_ID_OUT(fresh_wire_1800));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__99__DOLLAR__740$aRed(.PORT_ID_IN(fresh_wire_1801),
.PORT_ID_OUT(fresh_wire_1802));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__99__DOLLAR__740$andOps(.PORT_ID_IN0(fresh_wire_1803),
.PORT_ID_IN1(fresh_wire_1804),
.PORT_ID_OUT(fresh_wire_1805));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__99__DOLLAR__740$bRed(.PORT_ID_IN(fresh_wire_1806),
.PORT_ID_OUT(fresh_wire_1807));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__99__DOLLAR__742$aRed(.PORT_ID_IN(fresh_wire_1808),
.PORT_ID_OUT(fresh_wire_1809));

	CELL_TYPE_AND #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__99__DOLLAR__742$andOps(.PORT_ID_IN0(fresh_wire_1810),
.PORT_ID_IN1(fresh_wire_1811),
.PORT_ID_OUT(fresh_wire_1812));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_and__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__99__DOLLAR__742$bRed(.PORT_ID_IN(fresh_wire_1813),
.PORT_ID_OUT(fresh_wire_1814));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_or__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__124__DOLLAR__774$aRed(.PORT_ID_IN(fresh_wire_1815),
.PORT_ID_OUT(fresh_wire_1816));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_or__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__124__DOLLAR__774$bRed(.PORT_ID_IN(fresh_wire_1817),
.PORT_ID_OUT(fresh_wire_1818));

	CELL_TYPE_OR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_or__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__124__DOLLAR__774$orOps(.PORT_ID_IN0(fresh_wire_1819),
.PORT_ID_IN1(fresh_wire_1820),
.PORT_ID_OUT(fresh_wire_1821));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_or__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__126__DOLLAR__779$aRed(.PORT_ID_IN(fresh_wire_1822),
.PORT_ID_OUT(fresh_wire_1823));

	CELL_TYPE_ORR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_or__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__126__DOLLAR__779$bRed(.PORT_ID_IN(fresh_wire_1824),
.PORT_ID_OUT(fresh_wire_1825));

	CELL_TYPE_OR #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__logic_or__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__126__DOLLAR__779$orOps(.PORT_ID_IN0(fresh_wire_1826),
.PORT_ID_IN1(fresh_wire_1827),
.PORT_ID_OUT(fresh_wire_1828));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h1),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(2'h0),
.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__procdff__DOLLAR__3701$reg0(.PORT_ID_ARST(fresh_wire_1832),
.PORT_ID_CLK(fresh_wire_1831),
.PORT_ID_IN(fresh_wire_1829),
.PORT_ID_OUT(fresh_wire_1830));

	CELL_TYPE_REG #(.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(48'hxxxxxxxxxxxx),
.PARAM_WIDTH(32'h00000030)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__procdff__DOLLAR__3702$reg0(.PORT_ID_CLK(fresh_wire_1835),
.PORT_ID_IN(fresh_wire_1833),
.PORT_ID_OUT(fresh_wire_1834));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2382$mux0(.PORT_ID_IN0(fresh_wire_1836),
.PORT_ID_IN1(fresh_wire_1837),
.PORT_ID_OUT(fresh_wire_1838),
.PORT_ID_SEL(fresh_wire_1839));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2385$mux0(.PORT_ID_IN0(fresh_wire_1840),
.PORT_ID_IN1(fresh_wire_1841),
.PORT_ID_OUT(fresh_wire_1842),
.PORT_ID_SEL(fresh_wire_1843));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2388$mux0(.PORT_ID_IN0(fresh_wire_1844),
.PORT_ID_IN1(fresh_wire_1845),
.PORT_ID_OUT(fresh_wire_1846),
.PORT_ID_SEL(fresh_wire_1847));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2390$mux0(.PORT_ID_IN0(fresh_wire_1848),
.PORT_ID_IN1(fresh_wire_1849),
.PORT_ID_OUT(fresh_wire_1850),
.PORT_ID_SEL(fresh_wire_1851));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2393$mux0(.PORT_ID_IN0(fresh_wire_1852),
.PORT_ID_IN1(fresh_wire_1853),
.PORT_ID_OUT(fresh_wire_1854),
.PORT_ID_SEL(fresh_wire_1855));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2396$mux0(.PORT_ID_IN0(fresh_wire_1856),
.PORT_ID_IN1(fresh_wire_1857),
.PORT_ID_OUT(fresh_wire_1858),
.PORT_ID_SEL(fresh_wire_1859));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2399$mux0(.PORT_ID_IN0(fresh_wire_1860),
.PORT_ID_IN1(fresh_wire_1861),
.PORT_ID_OUT(fresh_wire_1862),
.PORT_ID_SEL(fresh_wire_1863));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2402$mux0(.PORT_ID_IN0(fresh_wire_1864),
.PORT_ID_IN1(fresh_wire_1865),
.PORT_ID_OUT(fresh_wire_1866),
.PORT_ID_SEL(fresh_wire_1867));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2406$mux0(.PORT_ID_IN0(fresh_wire_1868),
.PORT_ID_IN1(fresh_wire_1869),
.PORT_ID_OUT(fresh_wire_1870),
.PORT_ID_SEL(fresh_wire_1871));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2409$mux0(.PORT_ID_IN0(fresh_wire_1872),
.PORT_ID_IN1(fresh_wire_1873),
.PORT_ID_OUT(fresh_wire_1874),
.PORT_ID_SEL(fresh_wire_1875));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2412$mux0(.PORT_ID_IN0(fresh_wire_1876),
.PORT_ID_IN1(fresh_wire_1877),
.PORT_ID_OUT(fresh_wire_1878),
.PORT_ID_SEL(fresh_wire_1879));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2415$mux0(.PORT_ID_IN0(fresh_wire_1880),
.PORT_ID_IN1(fresh_wire_1881),
.PORT_ID_OUT(fresh_wire_1882),
.PORT_ID_SEL(fresh_wire_1883));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2418$mux0(.PORT_ID_IN0(fresh_wire_1884),
.PORT_ID_IN1(fresh_wire_1885),
.PORT_ID_OUT(fresh_wire_1886),
.PORT_ID_SEL(fresh_wire_1887));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000030)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2427$mux0(.PORT_ID_IN0(fresh_wire_1888),
.PORT_ID_IN1(fresh_wire_1889),
.PORT_ID_OUT(fresh_wire_1890),
.PORT_ID_SEL(fresh_wire_1891));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000030)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__procmux__DOLLAR__2430$mux0(.PORT_ID_IN0(fresh_wire_1892),
.PORT_ID_IN1(fresh_wire_1893),
.PORT_ID_OUT(fresh_wire_1894),
.PORT_ID_SEL(fresh_wire_1895));

	CELL_TYPE_SUB #(.PARAM_WIDTH(32'h00000002)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__sub__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__100__DOLLAR__743$op0(.PORT_ID_IN0(fresh_wire_1896),
.PORT_ID_IN1(fresh_wire_1897),
.PORT_ID_OUT(fresh_wire_1898));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$linebuffer_control$output_sr$__DOLLAR__sub__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__output_sr_unq1__DOT__v__COLON__100__DOLLAR__743__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(.PORT_ID_OUT(fresh_wire_1899));

	CELL_TYPE_NOT #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$__DOLLAR__not__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__mem_unq1__DOT__v__COLON__65__DOLLAR__575$op0(.PORT_ID_IN(fresh_wire_1900),
.PORT_ID_OUT(fresh_wire_1901));

	CELL_TYPE_NOT #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$__DOLLAR__not__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__mem_unq1__DOT__v__COLON__66__DOLLAR__576$op0(.PORT_ID_IN(fresh_wire_1902),
.PORT_ID_OUT(fresh_wire_1903));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__sram_512w_16b__DOT__v__COLON__38__DOLLAR__1114$op0(.PORT_ID_IN0(fresh_wire_1904),
.PORT_ID_IN1(fresh_wire_1905),
.PORT_ID_OUT(fresh_wire_1906));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__sram_512w_16b__DOT__v__COLON__40__DOLLAR__1116$op0(.PORT_ID_IN0(fresh_wire_1907),
.PORT_ID_IN1(fresh_wire_1908),
.PORT_ID_OUT(fresh_wire_1909));

	CELL_TYPE_REG #(.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(16'hxxxx),
.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procdff__DOLLAR__3630$reg0(.PORT_ID_CLK(fresh_wire_1912),
.PORT_ID_IN(fresh_wire_1910),
.PORT_ID_OUT(fresh_wire_1911));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1557$mux0(.PORT_ID_IN0(fresh_wire_1913),
.PORT_ID_IN1(fresh_wire_1914),
.PORT_ID_OUT(fresh_wire_1915),
.PORT_ID_SEL(fresh_wire_1916));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1567$mux0(.PORT_ID_IN0(fresh_wire_1917),
.PORT_ID_IN1(fresh_wire_1918),
.PORT_ID_OUT(fresh_wire_1919),
.PORT_ID_SEL(fresh_wire_1920));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1567__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(.PORT_ID_OUT(fresh_wire_1921));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1569$mux0(.PORT_ID_IN0(fresh_wire_1922),
.PORT_ID_IN1(fresh_wire_1923),
.PORT_ID_OUT(fresh_wire_1924),
.PORT_ID_SEL(fresh_wire_1925));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576$mux0(.PORT_ID_IN0(fresh_wire_1926),
.PORT_ID_IN1(fresh_wire_1927),
.PORT_ID_OUT(fresh_wire_1928),
.PORT_ID_SEL(fresh_wire_1929));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0$uConst(.PORT_ID_OUT(fresh_wire_1930));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10$uConst(.PORT_ID_OUT(fresh_wire_1931));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11$uConst(.PORT_ID_OUT(fresh_wire_1932));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12$uConst(.PORT_ID_OUT(fresh_wire_1933));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13$uConst(.PORT_ID_OUT(fresh_wire_1934));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14$uConst(.PORT_ID_OUT(fresh_wire_1935));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15$uConst(.PORT_ID_OUT(fresh_wire_1936));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1$uConst(.PORT_ID_OUT(fresh_wire_1937));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2$uConst(.PORT_ID_OUT(fresh_wire_1938));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3$uConst(.PORT_ID_OUT(fresh_wire_1939));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4$uConst(.PORT_ID_OUT(fresh_wire_1940));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5$uConst(.PORT_ID_OUT(fresh_wire_1941));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6$uConst(.PORT_ID_OUT(fresh_wire_1942));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7$uConst(.PORT_ID_OUT(fresh_wire_1943));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8$uConst(.PORT_ID_OUT(fresh_wire_1944));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9$uConst(.PORT_ID_OUT(fresh_wire_1945));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578$mux0(.PORT_ID_IN0(fresh_wire_1946),
.PORT_ID_IN1(fresh_wire_1947),
.PORT_ID_OUT(fresh_wire_1948),
.PORT_ID_SEL(fresh_wire_1949));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0$uConst(.PORT_ID_OUT(fresh_wire_1950));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10$uConst(.PORT_ID_OUT(fresh_wire_1951));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11$uConst(.PORT_ID_OUT(fresh_wire_1952));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12$uConst(.PORT_ID_OUT(fresh_wire_1953));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13$uConst(.PORT_ID_OUT(fresh_wire_1954));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14$uConst(.PORT_ID_OUT(fresh_wire_1955));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15$uConst(.PORT_ID_OUT(fresh_wire_1956));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1$uConst(.PORT_ID_OUT(fresh_wire_1957));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2$uConst(.PORT_ID_OUT(fresh_wire_1958));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3$uConst(.PORT_ID_OUT(fresh_wire_1959));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4$uConst(.PORT_ID_OUT(fresh_wire_1960));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5$uConst(.PORT_ID_OUT(fresh_wire_1961));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6$uConst(.PORT_ID_OUT(fresh_wire_1962));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7$uConst(.PORT_ID_OUT(fresh_wire_1963));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8$uConst(.PORT_ID_OUT(fresh_wire_1964));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9$uConst(.PORT_ID_OUT(fresh_wire_1965));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000009)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585$mux0(.PORT_ID_IN0(fresh_wire_1966),
.PORT_ID_IN1(fresh_wire_1967),
.PORT_ID_OUT(fresh_wire_1968),
.PORT_ID_SEL(fresh_wire_1969));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0$uConst(.PORT_ID_OUT(fresh_wire_1970));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1$uConst(.PORT_ID_OUT(fresh_wire_1971));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2$uConst(.PORT_ID_OUT(fresh_wire_1972));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3$uConst(.PORT_ID_OUT(fresh_wire_1973));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4$uConst(.PORT_ID_OUT(fresh_wire_1974));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5$uConst(.PORT_ID_OUT(fresh_wire_1975));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6$uConst(.PORT_ID_OUT(fresh_wire_1976));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7$uConst(.PORT_ID_OUT(fresh_wire_1977));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8$uConst(.PORT_ID_OUT(fresh_wire_1978));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000009)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587$mux0(.PORT_ID_IN0(fresh_wire_1979),
.PORT_ID_IN1(fresh_wire_1980),
.PORT_ID_OUT(fresh_wire_1981),
.PORT_ID_SEL(fresh_wire_1982));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0$uConst(.PORT_ID_OUT(fresh_wire_1983));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1$uConst(.PORT_ID_OUT(fresh_wire_1984));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2$uConst(.PORT_ID_OUT(fresh_wire_1985));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3$uConst(.PORT_ID_OUT(fresh_wire_1986));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4$uConst(.PORT_ID_OUT(fresh_wire_1987));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5$uConst(.PORT_ID_OUT(fresh_wire_1988));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6$uConst(.PORT_ID_OUT(fresh_wire_1989));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7$uConst(.PORT_ID_OUT(fresh_wire_1990));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst0$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8$uConst(.PORT_ID_OUT(fresh_wire_1991));

	CELL_TYPE_MEM #(.PARAM_HAS_INIT(1'h0),
.PARAM_MEM_DEPTH(32'h00000200),
.PARAM_MEM_WIDTH(32'h00000010)) mem_0x39$memory_core$mem_inst0$mem_inst$data_array$mem(.PORT_ID_CLK(fresh_wire_1992),
.PORT_ID_RADDR(fresh_wire_1993),
.PORT_ID_RDATA(fresh_wire_1994),
.PORT_ID_WADDR(fresh_wire_1995),
.PORT_ID_WDATA(fresh_wire_1996),
.PORT_ID_WEN(fresh_wire_1997));

	CELL_TYPE_NOT #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$__DOLLAR__not__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__mem_unq1__DOT__v__COLON__65__DOLLAR__575$op0(.PORT_ID_IN(fresh_wire_1998),
.PORT_ID_OUT(fresh_wire_1999));

	CELL_TYPE_NOT #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$__DOLLAR__not__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__mem_unq1__DOT__v__COLON__66__DOLLAR__576$op0(.PORT_ID_IN(fresh_wire_2000),
.PORT_ID_OUT(fresh_wire_2001));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__sram_512w_16b__DOT__v__COLON__38__DOLLAR__1114$op0(.PORT_ID_IN0(fresh_wire_2002),
.PORT_ID_IN1(fresh_wire_2003),
.PORT_ID_OUT(fresh_wire_2004));

	CELL_TYPE_EQ #(.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__eq__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__sram_512w_16b__DOT__v__COLON__40__DOLLAR__1116$op0(.PORT_ID_IN0(fresh_wire_2005),
.PORT_ID_IN1(fresh_wire_2006),
.PORT_ID_OUT(fresh_wire_2007));

	CELL_TYPE_REG #(.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(16'hxxxx),
.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procdff__DOLLAR__3630$reg0(.PORT_ID_CLK(fresh_wire_2010),
.PORT_ID_IN(fresh_wire_2008),
.PORT_ID_OUT(fresh_wire_2009));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1557$mux0(.PORT_ID_IN0(fresh_wire_2011),
.PORT_ID_IN1(fresh_wire_2012),
.PORT_ID_OUT(fresh_wire_2013),
.PORT_ID_SEL(fresh_wire_2014));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1567$mux0(.PORT_ID_IN0(fresh_wire_2015),
.PORT_ID_IN1(fresh_wire_2016),
.PORT_ID_OUT(fresh_wire_2017),
.PORT_ID_SEL(fresh_wire_2018));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1567__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(.PORT_ID_OUT(fresh_wire_2019));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1569$mux0(.PORT_ID_IN0(fresh_wire_2020),
.PORT_ID_IN1(fresh_wire_2021),
.PORT_ID_OUT(fresh_wire_2022),
.PORT_ID_SEL(fresh_wire_2023));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576$mux0(.PORT_ID_IN0(fresh_wire_2024),
.PORT_ID_IN1(fresh_wire_2025),
.PORT_ID_OUT(fresh_wire_2026),
.PORT_ID_SEL(fresh_wire_2027));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0$uConst(.PORT_ID_OUT(fresh_wire_2028));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10$uConst(.PORT_ID_OUT(fresh_wire_2029));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11$uConst(.PORT_ID_OUT(fresh_wire_2030));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12$uConst(.PORT_ID_OUT(fresh_wire_2031));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13$uConst(.PORT_ID_OUT(fresh_wire_2032));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14$uConst(.PORT_ID_OUT(fresh_wire_2033));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15$uConst(.PORT_ID_OUT(fresh_wire_2034));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1$uConst(.PORT_ID_OUT(fresh_wire_2035));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2$uConst(.PORT_ID_OUT(fresh_wire_2036));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3$uConst(.PORT_ID_OUT(fresh_wire_2037));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4$uConst(.PORT_ID_OUT(fresh_wire_2038));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5$uConst(.PORT_ID_OUT(fresh_wire_2039));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6$uConst(.PORT_ID_OUT(fresh_wire_2040));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7$uConst(.PORT_ID_OUT(fresh_wire_2041));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8$uConst(.PORT_ID_OUT(fresh_wire_2042));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1576__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9$uConst(.PORT_ID_OUT(fresh_wire_2043));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000010)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578$mux0(.PORT_ID_IN0(fresh_wire_2044),
.PORT_ID_IN1(fresh_wire_2045),
.PORT_ID_OUT(fresh_wire_2046),
.PORT_ID_SEL(fresh_wire_2047));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0$uConst(.PORT_ID_OUT(fresh_wire_2048));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10$uConst(.PORT_ID_OUT(fresh_wire_2049));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11$uConst(.PORT_ID_OUT(fresh_wire_2050));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12$uConst(.PORT_ID_OUT(fresh_wire_2051));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13$uConst(.PORT_ID_OUT(fresh_wire_2052));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14$uConst(.PORT_ID_OUT(fresh_wire_2053));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15$uConst(.PORT_ID_OUT(fresh_wire_2054));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1$uConst(.PORT_ID_OUT(fresh_wire_2055));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2$uConst(.PORT_ID_OUT(fresh_wire_2056));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3$uConst(.PORT_ID_OUT(fresh_wire_2057));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4$uConst(.PORT_ID_OUT(fresh_wire_2058));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5$uConst(.PORT_ID_OUT(fresh_wire_2059));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6$uConst(.PORT_ID_OUT(fresh_wire_2060));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7$uConst(.PORT_ID_OUT(fresh_wire_2061));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8$uConst(.PORT_ID_OUT(fresh_wire_2062));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1578__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9$uConst(.PORT_ID_OUT(fresh_wire_2063));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000009)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585$mux0(.PORT_ID_IN0(fresh_wire_2064),
.PORT_ID_IN1(fresh_wire_2065),
.PORT_ID_OUT(fresh_wire_2066),
.PORT_ID_SEL(fresh_wire_2067));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0$uConst(.PORT_ID_OUT(fresh_wire_2068));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1$uConst(.PORT_ID_OUT(fresh_wire_2069));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2$uConst(.PORT_ID_OUT(fresh_wire_2070));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3$uConst(.PORT_ID_OUT(fresh_wire_2071));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4$uConst(.PORT_ID_OUT(fresh_wire_2072));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5$uConst(.PORT_ID_OUT(fresh_wire_2073));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6$uConst(.PORT_ID_OUT(fresh_wire_2074));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7$uConst(.PORT_ID_OUT(fresh_wire_2075));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1585__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8$uConst(.PORT_ID_OUT(fresh_wire_2076));

	CELL_TYPE_MUX #(.PARAM_WIDTH(32'h00000009)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587$mux0(.PORT_ID_IN0(fresh_wire_2077),
.PORT_ID_IN1(fresh_wire_2078),
.PORT_ID_OUT(fresh_wire_2079),
.PORT_ID_SEL(fresh_wire_2080));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0$uConst(.PORT_ID_OUT(fresh_wire_2081));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1$uConst(.PORT_ID_OUT(fresh_wire_2082));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2$uConst(.PORT_ID_OUT(fresh_wire_2083));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3$uConst(.PORT_ID_OUT(fresh_wire_2084));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4$uConst(.PORT_ID_OUT(fresh_wire_2085));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5$uConst(.PORT_ID_OUT(fresh_wire_2086));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6$uConst(.PORT_ID_OUT(fresh_wire_2087));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7$uConst(.PORT_ID_OUT(fresh_wire_2088));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'hx),
.PARAM_WIDTH(32'h00000001)) mem_0x39$memory_core$mem_inst1$mem_inst$__DOLLAR__procmux__DOLLAR__1587__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8$uConst(.PORT_ID_OUT(fresh_wire_2089));

	CELL_TYPE_MEM #(.PARAM_HAS_INIT(1'h0),
.PARAM_MEM_DEPTH(32'h00000200),
.PARAM_MEM_WIDTH(32'h00000010)) mem_0x39$memory_core$mem_inst1$mem_inst$data_array$mem(.PORT_ID_CLK(fresh_wire_2090),
.PORT_ID_RADDR(fresh_wire_2091),
.PORT_ID_RDATA(fresh_wire_2092),
.PORT_ID_WADDR(fresh_wire_2093),
.PORT_ID_WDATA(fresh_wire_2094),
.PORT_ID_WEN(fresh_wire_2095));

	CELL_TYPE_REG #(.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(16'hxxxx),
.PARAM_WIDTH(32'h00000010)) mem_0x39$sb_inst_busBUS16_row0$__DOLLAR__procdff__DOLLAR__3697$reg0(.PORT_ID_CLK(fresh_wire_2098),
.PORT_ID_IN(fresh_wire_2096),
.PORT_ID_OUT(fresh_wire_2097));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T0_in_port_cell(.PORT_ID_IN(pad_S0_T0_in),
.PORT_ID_OUT(fresh_wire_20));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T0_out_port_cell(.PORT_ID_IN(fresh_wire_21),
.PORT_ID_OUT(pad_S0_T0_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T10_in_port_cell(.PORT_ID_IN(pad_S0_T10_in),
.PORT_ID_OUT(fresh_wire_22));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T10_out_port_cell(.PORT_ID_IN(fresh_wire_23),
.PORT_ID_OUT(pad_S0_T10_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T11_in_port_cell(.PORT_ID_IN(pad_S0_T11_in),
.PORT_ID_OUT(fresh_wire_24));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T11_out_port_cell(.PORT_ID_IN(fresh_wire_25),
.PORT_ID_OUT(pad_S0_T11_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T12_in_port_cell(.PORT_ID_IN(pad_S0_T12_in),
.PORT_ID_OUT(fresh_wire_26));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T12_out_port_cell(.PORT_ID_IN(fresh_wire_27),
.PORT_ID_OUT(pad_S0_T12_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T13_in_port_cell(.PORT_ID_IN(pad_S0_T13_in),
.PORT_ID_OUT(fresh_wire_28));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T13_out_port_cell(.PORT_ID_IN(fresh_wire_29),
.PORT_ID_OUT(pad_S0_T13_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T14_in_port_cell(.PORT_ID_IN(pad_S0_T14_in),
.PORT_ID_OUT(fresh_wire_30));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T14_out_port_cell(.PORT_ID_IN(fresh_wire_31),
.PORT_ID_OUT(pad_S0_T14_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T15_in_port_cell(.PORT_ID_IN(pad_S0_T15_in),
.PORT_ID_OUT(fresh_wire_32));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T15_out_port_cell(.PORT_ID_IN(fresh_wire_33),
.PORT_ID_OUT(pad_S0_T15_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T1_in_port_cell(.PORT_ID_IN(pad_S0_T1_in),
.PORT_ID_OUT(fresh_wire_34));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T1_out_port_cell(.PORT_ID_IN(fresh_wire_35),
.PORT_ID_OUT(pad_S0_T1_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T2_in_port_cell(.PORT_ID_IN(pad_S0_T2_in),
.PORT_ID_OUT(fresh_wire_36));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T2_out_port_cell(.PORT_ID_IN(fresh_wire_37),
.PORT_ID_OUT(pad_S0_T2_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T3_in_port_cell(.PORT_ID_IN(pad_S0_T3_in),
.PORT_ID_OUT(fresh_wire_38));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T3_out_port_cell(.PORT_ID_IN(fresh_wire_39),
.PORT_ID_OUT(pad_S0_T3_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T4_in_port_cell(.PORT_ID_IN(pad_S0_T4_in),
.PORT_ID_OUT(fresh_wire_40));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T4_out_port_cell(.PORT_ID_IN(fresh_wire_41),
.PORT_ID_OUT(pad_S0_T4_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T5_in_port_cell(.PORT_ID_IN(pad_S0_T5_in),
.PORT_ID_OUT(fresh_wire_42));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T5_out_port_cell(.PORT_ID_IN(fresh_wire_43),
.PORT_ID_OUT(pad_S0_T5_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T6_in_port_cell(.PORT_ID_IN(pad_S0_T6_in),
.PORT_ID_OUT(fresh_wire_44));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T6_out_port_cell(.PORT_ID_IN(fresh_wire_45),
.PORT_ID_OUT(pad_S0_T6_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T7_in_port_cell(.PORT_ID_IN(pad_S0_T7_in),
.PORT_ID_OUT(fresh_wire_46));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T7_out_port_cell(.PORT_ID_IN(fresh_wire_47),
.PORT_ID_OUT(pad_S0_T7_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T8_in_port_cell(.PORT_ID_IN(pad_S0_T8_in),
.PORT_ID_OUT(fresh_wire_48));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T8_out_port_cell(.PORT_ID_IN(fresh_wire_49),
.PORT_ID_OUT(pad_S0_T8_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T9_in_port_cell(.PORT_ID_IN(pad_S0_T9_in),
.PORT_ID_OUT(fresh_wire_50));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T9_out_port_cell(.PORT_ID_IN(fresh_wire_51),
.PORT_ID_OUT(pad_S0_T9_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T0_in_port_cell(.PORT_ID_IN(pad_S1_T0_in),
.PORT_ID_OUT(fresh_wire_52));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T0_out_port_cell(.PORT_ID_IN(fresh_wire_53),
.PORT_ID_OUT(pad_S1_T0_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T10_in_port_cell(.PORT_ID_IN(pad_S1_T10_in),
.PORT_ID_OUT(fresh_wire_54));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T10_out_port_cell(.PORT_ID_IN(fresh_wire_55),
.PORT_ID_OUT(pad_S1_T10_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T11_in_port_cell(.PORT_ID_IN(pad_S1_T11_in),
.PORT_ID_OUT(fresh_wire_56));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T11_out_port_cell(.PORT_ID_IN(fresh_wire_57),
.PORT_ID_OUT(pad_S1_T11_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T12_in_port_cell(.PORT_ID_IN(pad_S1_T12_in),
.PORT_ID_OUT(fresh_wire_58));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T12_out_port_cell(.PORT_ID_IN(fresh_wire_59),
.PORT_ID_OUT(pad_S1_T12_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T13_in_port_cell(.PORT_ID_IN(pad_S1_T13_in),
.PORT_ID_OUT(fresh_wire_60));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T13_out_port_cell(.PORT_ID_IN(fresh_wire_61),
.PORT_ID_OUT(pad_S1_T13_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T14_in_port_cell(.PORT_ID_IN(pad_S1_T14_in),
.PORT_ID_OUT(fresh_wire_62));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T14_out_port_cell(.PORT_ID_IN(fresh_wire_63),
.PORT_ID_OUT(pad_S1_T14_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T15_in_port_cell(.PORT_ID_IN(pad_S1_T15_in),
.PORT_ID_OUT(fresh_wire_64));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T15_out_port_cell(.PORT_ID_IN(fresh_wire_65),
.PORT_ID_OUT(pad_S1_T15_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T1_in_port_cell(.PORT_ID_IN(pad_S1_T1_in),
.PORT_ID_OUT(fresh_wire_66));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T1_out_port_cell(.PORT_ID_IN(fresh_wire_67),
.PORT_ID_OUT(pad_S1_T1_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T2_in_port_cell(.PORT_ID_IN(pad_S1_T2_in),
.PORT_ID_OUT(fresh_wire_68));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T2_out_port_cell(.PORT_ID_IN(fresh_wire_69),
.PORT_ID_OUT(pad_S1_T2_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T3_in_port_cell(.PORT_ID_IN(pad_S1_T3_in),
.PORT_ID_OUT(fresh_wire_70));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T3_out_port_cell(.PORT_ID_IN(fresh_wire_71),
.PORT_ID_OUT(pad_S1_T3_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T4_in_port_cell(.PORT_ID_IN(pad_S1_T4_in),
.PORT_ID_OUT(fresh_wire_72));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T4_out_port_cell(.PORT_ID_IN(fresh_wire_73),
.PORT_ID_OUT(pad_S1_T4_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T5_in_port_cell(.PORT_ID_IN(pad_S1_T5_in),
.PORT_ID_OUT(fresh_wire_74));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T5_out_port_cell(.PORT_ID_IN(fresh_wire_75),
.PORT_ID_OUT(pad_S1_T5_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T6_in_port_cell(.PORT_ID_IN(pad_S1_T6_in),
.PORT_ID_OUT(fresh_wire_76));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T6_out_port_cell(.PORT_ID_IN(fresh_wire_77),
.PORT_ID_OUT(pad_S1_T6_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T7_in_port_cell(.PORT_ID_IN(pad_S1_T7_in),
.PORT_ID_OUT(fresh_wire_78));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T7_out_port_cell(.PORT_ID_IN(fresh_wire_79),
.PORT_ID_OUT(pad_S1_T7_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T8_in_port_cell(.PORT_ID_IN(pad_S1_T8_in),
.PORT_ID_OUT(fresh_wire_80));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T8_out_port_cell(.PORT_ID_IN(fresh_wire_81),
.PORT_ID_OUT(pad_S1_T8_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T9_in_port_cell(.PORT_ID_IN(pad_S1_T9_in),
.PORT_ID_OUT(fresh_wire_82));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T9_out_port_cell(.PORT_ID_IN(fresh_wire_83),
.PORT_ID_OUT(pad_S1_T9_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T0_in_port_cell(.PORT_ID_IN(pad_S2_T0_in),
.PORT_ID_OUT(fresh_wire_84));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T0_out_port_cell(.PORT_ID_IN(fresh_wire_85),
.PORT_ID_OUT(pad_S2_T0_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T10_in_port_cell(.PORT_ID_IN(pad_S2_T10_in),
.PORT_ID_OUT(fresh_wire_86));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T10_out_port_cell(.PORT_ID_IN(fresh_wire_87),
.PORT_ID_OUT(pad_S2_T10_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T11_in_port_cell(.PORT_ID_IN(pad_S2_T11_in),
.PORT_ID_OUT(fresh_wire_88));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T11_out_port_cell(.PORT_ID_IN(fresh_wire_89),
.PORT_ID_OUT(pad_S2_T11_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T12_in_port_cell(.PORT_ID_IN(pad_S2_T12_in),
.PORT_ID_OUT(fresh_wire_90));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T12_out_port_cell(.PORT_ID_IN(fresh_wire_91),
.PORT_ID_OUT(pad_S2_T12_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T13_in_port_cell(.PORT_ID_IN(pad_S2_T13_in),
.PORT_ID_OUT(fresh_wire_92));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T13_out_port_cell(.PORT_ID_IN(fresh_wire_93),
.PORT_ID_OUT(pad_S2_T13_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T14_in_port_cell(.PORT_ID_IN(pad_S2_T14_in),
.PORT_ID_OUT(fresh_wire_94));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T14_out_port_cell(.PORT_ID_IN(fresh_wire_95),
.PORT_ID_OUT(pad_S2_T14_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T15_in_port_cell(.PORT_ID_IN(pad_S2_T15_in),
.PORT_ID_OUT(fresh_wire_96));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T15_out_port_cell(.PORT_ID_IN(fresh_wire_97),
.PORT_ID_OUT(pad_S2_T15_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T1_in_port_cell(.PORT_ID_IN(pad_S2_T1_in),
.PORT_ID_OUT(fresh_wire_98));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T1_out_port_cell(.PORT_ID_IN(fresh_wire_99),
.PORT_ID_OUT(pad_S2_T1_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T2_in_port_cell(.PORT_ID_IN(pad_S2_T2_in),
.PORT_ID_OUT(fresh_wire_100));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T2_out_port_cell(.PORT_ID_IN(fresh_wire_101),
.PORT_ID_OUT(pad_S2_T2_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T3_in_port_cell(.PORT_ID_IN(pad_S2_T3_in),
.PORT_ID_OUT(fresh_wire_102));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T3_out_port_cell(.PORT_ID_IN(fresh_wire_103),
.PORT_ID_OUT(pad_S2_T3_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T4_in_port_cell(.PORT_ID_IN(pad_S2_T4_in),
.PORT_ID_OUT(fresh_wire_104));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T4_out_port_cell(.PORT_ID_IN(fresh_wire_105),
.PORT_ID_OUT(pad_S2_T4_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T5_in_port_cell(.PORT_ID_IN(pad_S2_T5_in),
.PORT_ID_OUT(fresh_wire_106));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T5_out_port_cell(.PORT_ID_IN(fresh_wire_107),
.PORT_ID_OUT(pad_S2_T5_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T6_in_port_cell(.PORT_ID_IN(pad_S2_T6_in),
.PORT_ID_OUT(fresh_wire_108));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T6_out_port_cell(.PORT_ID_IN(fresh_wire_109),
.PORT_ID_OUT(pad_S2_T6_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T7_in_port_cell(.PORT_ID_IN(pad_S2_T7_in),
.PORT_ID_OUT(fresh_wire_110));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T7_out_port_cell(.PORT_ID_IN(fresh_wire_111),
.PORT_ID_OUT(pad_S2_T7_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T8_in_port_cell(.PORT_ID_IN(pad_S2_T8_in),
.PORT_ID_OUT(fresh_wire_112));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T8_out_port_cell(.PORT_ID_IN(fresh_wire_113),
.PORT_ID_OUT(pad_S2_T8_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T9_in_port_cell(.PORT_ID_IN(pad_S2_T9_in),
.PORT_ID_OUT(fresh_wire_114));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T9_out_port_cell(.PORT_ID_IN(fresh_wire_115),
.PORT_ID_OUT(pad_S2_T9_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T0_in_port_cell(.PORT_ID_IN(pad_S3_T0_in),
.PORT_ID_OUT(fresh_wire_116));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T0_out_port_cell(.PORT_ID_IN(fresh_wire_117),
.PORT_ID_OUT(pad_S3_T0_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T10_in_port_cell(.PORT_ID_IN(pad_S3_T10_in),
.PORT_ID_OUT(fresh_wire_118));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T10_out_port_cell(.PORT_ID_IN(fresh_wire_119),
.PORT_ID_OUT(pad_S3_T10_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T11_in_port_cell(.PORT_ID_IN(pad_S3_T11_in),
.PORT_ID_OUT(fresh_wire_120));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T11_out_port_cell(.PORT_ID_IN(fresh_wire_121),
.PORT_ID_OUT(pad_S3_T11_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T12_in_port_cell(.PORT_ID_IN(pad_S3_T12_in),
.PORT_ID_OUT(fresh_wire_122));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T12_out_port_cell(.PORT_ID_IN(fresh_wire_123),
.PORT_ID_OUT(pad_S3_T12_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T13_in_port_cell(.PORT_ID_IN(pad_S3_T13_in),
.PORT_ID_OUT(fresh_wire_124));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T13_out_port_cell(.PORT_ID_IN(fresh_wire_125),
.PORT_ID_OUT(pad_S3_T13_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T14_in_port_cell(.PORT_ID_IN(pad_S3_T14_in),
.PORT_ID_OUT(fresh_wire_126));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T14_out_port_cell(.PORT_ID_IN(fresh_wire_127),
.PORT_ID_OUT(pad_S3_T14_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T15_in_port_cell(.PORT_ID_IN(pad_S3_T15_in),
.PORT_ID_OUT(fresh_wire_128));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T15_out_port_cell(.PORT_ID_IN(fresh_wire_129),
.PORT_ID_OUT(pad_S3_T15_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T1_in_port_cell(.PORT_ID_IN(pad_S3_T1_in),
.PORT_ID_OUT(fresh_wire_130));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T1_out_port_cell(.PORT_ID_IN(fresh_wire_131),
.PORT_ID_OUT(pad_S3_T1_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T2_in_port_cell(.PORT_ID_IN(pad_S3_T2_in),
.PORT_ID_OUT(fresh_wire_132));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T2_out_port_cell(.PORT_ID_IN(fresh_wire_133),
.PORT_ID_OUT(pad_S3_T2_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T3_in_port_cell(.PORT_ID_IN(pad_S3_T3_in),
.PORT_ID_OUT(fresh_wire_134));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T3_out_port_cell(.PORT_ID_IN(fresh_wire_135),
.PORT_ID_OUT(pad_S3_T3_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T4_in_port_cell(.PORT_ID_IN(pad_S3_T4_in),
.PORT_ID_OUT(fresh_wire_136));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T4_out_port_cell(.PORT_ID_IN(fresh_wire_137),
.PORT_ID_OUT(pad_S3_T4_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T5_in_port_cell(.PORT_ID_IN(pad_S3_T5_in),
.PORT_ID_OUT(fresh_wire_138));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T5_out_port_cell(.PORT_ID_IN(fresh_wire_139),
.PORT_ID_OUT(pad_S3_T5_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T6_in_port_cell(.PORT_ID_IN(pad_S3_T6_in),
.PORT_ID_OUT(fresh_wire_140));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T6_out_port_cell(.PORT_ID_IN(fresh_wire_141),
.PORT_ID_OUT(pad_S3_T6_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T7_in_port_cell(.PORT_ID_IN(pad_S3_T7_in),
.PORT_ID_OUT(fresh_wire_142));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T7_out_port_cell(.PORT_ID_IN(fresh_wire_143),
.PORT_ID_OUT(pad_S3_T7_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T8_in_port_cell(.PORT_ID_IN(pad_S3_T8_in),
.PORT_ID_OUT(fresh_wire_144));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T8_out_port_cell(.PORT_ID_IN(fresh_wire_145),
.PORT_ID_OUT(pad_S3_T8_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T9_in_port_cell(.PORT_ID_IN(pad_S3_T9_in),
.PORT_ID_OUT(fresh_wire_146));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T9_out_port_cell(.PORT_ID_IN(fresh_wire_147),
.PORT_ID_OUT(pad_S3_T9_out));

	CELL_TYPE_REG #(.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(16'hxxxx),
.PARAM_WIDTH(32'h00000010)) pe_0x15$sb_wide$__DOLLAR__procdff__DOLLAR__3692$reg0(.PORT_ID_CLK(fresh_wire_2101),
.PORT_ID_IN(fresh_wire_2099),
.PORT_ID_OUT(fresh_wire_2100));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000011),
.PARAM_OUT_WIDTH(32'h00000022)) pe_0x15$test_pe$test_pe_comp$test_mult_add$__DOLLAR__mul__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__1503$extendA(.PORT_ID_IN(fresh_wire_2102),
.PORT_ID_OUT(fresh_wire_2103));

	CELL_TYPE_MUL #(.PARAM_WIDTH(32'h00000022)) pe_0x15$test_pe$test_pe_comp$test_mult_add$__DOLLAR__mul__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__1503$op0(.PORT_ID_IN0(fresh_wire_2104),
.PORT_ID_IN1(fresh_wire_2105),
.PORT_ID_OUT(fresh_wire_2106));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000011),
.PARAM_OUT_WIDTH(32'h00000022)) pe_0x16$test_pe$test_pe_comp$test_mult_add$__DOLLAR__mul__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__1503$extendA(.PORT_ID_IN(fresh_wire_2107),
.PORT_ID_OUT(fresh_wire_2108));

	CELL_TYPE_MUL #(.PARAM_WIDTH(32'h00000022)) pe_0x16$test_pe$test_pe_comp$test_mult_add$__DOLLAR__mul__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__1503$op0(.PORT_ID_IN0(fresh_wire_2109),
.PORT_ID_IN1(fresh_wire_2110),
.PORT_ID_OUT(fresh_wire_2111));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000011),
.PARAM_OUT_WIDTH(32'h00000022)) pe_0x17$test_pe$test_pe_comp$test_mult_add$__DOLLAR__mul__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__1503$extendA(.PORT_ID_IN(fresh_wire_2112),
.PORT_ID_OUT(fresh_wire_2113));

	CELL_TYPE_MUL #(.PARAM_WIDTH(32'h00000022)) pe_0x17$test_pe$test_pe_comp$test_mult_add$__DOLLAR__mul__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__1503$op0(.PORT_ID_IN0(fresh_wire_2114),
.PORT_ID_IN1(fresh_wire_2115),
.PORT_ID_OUT(fresh_wire_2116));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) pe_0x19$test_pe$test_lut$self__DOT__res__DOLLAR__bit_const_0(.PORT_ID_OUT(fresh_wire_2117));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000011)) pe_0x28$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$extendA(.PORT_ID_IN(fresh_wire_2118),
.PORT_ID_OUT(fresh_wire_2119));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000011)) pe_0x28$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$extendB(.PORT_ID_IN(fresh_wire_2120),
.PORT_ID_OUT(fresh_wire_2121));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000011)) pe_0x28$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$op0(.PORT_ID_IN0(fresh_wire_2122),
.PORT_ID_IN1(fresh_wire_2123),
.PORT_ID_OUT(fresh_wire_2124));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000011)) pe_0x28$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1495$op0(.PORT_ID_IN0(fresh_wire_2125),
.PORT_ID_IN1(fresh_wire_2126),
.PORT_ID_OUT(fresh_wire_2127));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000011)) pe_0x29$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$extendA(.PORT_ID_IN(fresh_wire_2128),
.PORT_ID_OUT(fresh_wire_2129));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000011)) pe_0x29$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$extendB(.PORT_ID_IN(fresh_wire_2130),
.PORT_ID_OUT(fresh_wire_2131));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000011)) pe_0x29$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$op0(.PORT_ID_IN0(fresh_wire_2132),
.PORT_ID_IN1(fresh_wire_2133),
.PORT_ID_OUT(fresh_wire_2134));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000011)) pe_0x29$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1495$op0(.PORT_ID_IN0(fresh_wire_2135),
.PORT_ID_IN1(fresh_wire_2136),
.PORT_ID_OUT(fresh_wire_2137));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000011),
.PARAM_OUT_WIDTH(32'h00000022)) pe_0x2A$test_pe$test_pe_comp$test_mult_add$__DOLLAR__mul__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__1503$extendA(.PORT_ID_IN(fresh_wire_2138),
.PORT_ID_OUT(fresh_wire_2139));

	CELL_TYPE_MUL #(.PARAM_WIDTH(32'h00000022)) pe_0x2A$test_pe$test_pe_comp$test_mult_add$__DOLLAR__mul__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__1503$op0(.PORT_ID_IN0(fresh_wire_2140),
.PORT_ID_IN1(fresh_wire_2141),
.PORT_ID_OUT(fresh_wire_2142));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h0),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(16'h0000),
.PARAM_WIDTH(32'h00000010)) pe_0x2B$test_pe$test_opt_reg_a$__DOLLAR__procdff__DOLLAR__3625$reg0(.PORT_ID_ARST(fresh_wire_2146),
.PORT_ID_CLK(fresh_wire_2145),
.PORT_ID_IN(fresh_wire_2143),
.PORT_ID_OUT(fresh_wire_2144));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000011),
.PARAM_OUT_WIDTH(32'h00000022)) pe_0x2B$test_pe$test_pe_comp$test_mult_add$__DOLLAR__mul__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__1503$extendA(.PORT_ID_IN(fresh_wire_2147),
.PORT_ID_OUT(fresh_wire_2148));

	CELL_TYPE_MUL #(.PARAM_WIDTH(32'h00000022)) pe_0x2B$test_pe$test_pe_comp$test_mult_add$__DOLLAR__mul__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__1503$op0(.PORT_ID_IN0(fresh_wire_2149),
.PORT_ID_IN1(fresh_wire_2150),
.PORT_ID_OUT(fresh_wire_2151));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000011)) pe_0x36$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$extendA(.PORT_ID_IN(fresh_wire_2152),
.PORT_ID_OUT(fresh_wire_2153));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000011)) pe_0x36$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$extendB(.PORT_ID_IN(fresh_wire_2154),
.PORT_ID_OUT(fresh_wire_2155));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000011)) pe_0x36$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$op0(.PORT_ID_IN0(fresh_wire_2156),
.PORT_ID_IN1(fresh_wire_2157),
.PORT_ID_OUT(fresh_wire_2158));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000011)) pe_0x36$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1495$op0(.PORT_ID_IN0(fresh_wire_2159),
.PORT_ID_IN1(fresh_wire_2160),
.PORT_ID_OUT(fresh_wire_2161));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000011)) pe_0x37$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$extendA(.PORT_ID_IN(fresh_wire_2162),
.PORT_ID_OUT(fresh_wire_2163));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000011)) pe_0x37$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$extendB(.PORT_ID_IN(fresh_wire_2164),
.PORT_ID_OUT(fresh_wire_2165));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000011)) pe_0x37$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$op0(.PORT_ID_IN0(fresh_wire_2166),
.PORT_ID_IN1(fresh_wire_2167),
.PORT_ID_OUT(fresh_wire_2168));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000011)) pe_0x37$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1495$op0(.PORT_ID_IN0(fresh_wire_2169),
.PORT_ID_IN1(fresh_wire_2170),
.PORT_ID_OUT(fresh_wire_2171));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000011),
.PARAM_OUT_WIDTH(32'h00000022)) pe_0x38$test_pe$test_pe_comp$test_mult_add$__DOLLAR__mul__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__1503$extendA(.PORT_ID_IN(fresh_wire_2172),
.PORT_ID_OUT(fresh_wire_2173));

	CELL_TYPE_MUL #(.PARAM_WIDTH(32'h00000022)) pe_0x38$test_pe$test_pe_comp$test_mult_add$__DOLLAR__mul__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__1503$op0(.PORT_ID_IN0(fresh_wire_2174),
.PORT_ID_IN1(fresh_wire_2175),
.PORT_ID_OUT(fresh_wire_2176));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h1),
.PARAM_WIDTH(32'h00000001)) pe_0x3A$test_pe$test_lut$self__DOT__res__DOLLAR__bit_const_0(.PORT_ID_OUT(fresh_wire_2177));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000011)) pe_0x3B$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$extendA(.PORT_ID_IN(fresh_wire_2178),
.PORT_ID_OUT(fresh_wire_2179));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000011)) pe_0x3B$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$op0(.PORT_ID_IN0(fresh_wire_2180),
.PORT_ID_IN1(fresh_wire_2181),
.PORT_ID_OUT(fresh_wire_2182));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000011)) pe_0x3B$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1495$op0(.PORT_ID_IN0(fresh_wire_2183),
.PORT_ID_IN1(fresh_wire_2184),
.PORT_ID_OUT(fresh_wire_2185));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000011)) pe_0x48$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$extendA(.PORT_ID_IN(fresh_wire_2186),
.PORT_ID_OUT(fresh_wire_2187));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000011)) pe_0x48$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$extendB(.PORT_ID_IN(fresh_wire_2188),
.PORT_ID_OUT(fresh_wire_2189));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000011)) pe_0x48$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$op0(.PORT_ID_IN0(fresh_wire_2190),
.PORT_ID_IN1(fresh_wire_2191),
.PORT_ID_OUT(fresh_wire_2192));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000011)) pe_0x48$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1495$op0(.PORT_ID_IN0(fresh_wire_2193),
.PORT_ID_IN1(fresh_wire_2194),
.PORT_ID_OUT(fresh_wire_2195));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000011)) pe_0x49$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$extendA(.PORT_ID_IN(fresh_wire_2196),
.PORT_ID_OUT(fresh_wire_2197));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000011)) pe_0x49$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$extendB(.PORT_ID_IN(fresh_wire_2198),
.PORT_ID_OUT(fresh_wire_2199));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000011)) pe_0x49$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$op0(.PORT_ID_IN0(fresh_wire_2200),
.PORT_ID_IN1(fresh_wire_2201),
.PORT_ID_OUT(fresh_wire_2202));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000011)) pe_0x49$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1495$op0(.PORT_ID_IN0(fresh_wire_2203),
.PORT_ID_IN1(fresh_wire_2204),
.PORT_ID_OUT(fresh_wire_2205));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000011)) pe_0x4A$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$extendA(.PORT_ID_IN(fresh_wire_2206),
.PORT_ID_OUT(fresh_wire_2207));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000011)) pe_0x4A$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$extendB(.PORT_ID_IN(fresh_wire_2208),
.PORT_ID_OUT(fresh_wire_2209));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000011)) pe_0x4A$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$op0(.PORT_ID_IN0(fresh_wire_2210),
.PORT_ID_IN1(fresh_wire_2211),
.PORT_ID_OUT(fresh_wire_2212));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000011)) pe_0x4A$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1495$op0(.PORT_ID_IN0(fresh_wire_2213),
.PORT_ID_IN1(fresh_wire_2214),
.PORT_ID_OUT(fresh_wire_2215));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000011),
.PARAM_OUT_WIDTH(32'h00000022)) pe_0x4B$test_pe$test_pe_comp$test_mult_add$__DOLLAR__mul__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__1503$extendA(.PORT_ID_IN(fresh_wire_2216),
.PORT_ID_OUT(fresh_wire_2217));

	CELL_TYPE_MUL #(.PARAM_WIDTH(32'h00000022)) pe_0x4B$test_pe$test_pe_comp$test_mult_add$__DOLLAR__mul__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__1503$op0(.PORT_ID_IN0(fresh_wire_2218),
.PORT_ID_IN1(fresh_wire_2219),
.PORT_ID_OUT(fresh_wire_2220));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h0),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(16'h0000),
.PARAM_WIDTH(32'h00000010)) pe_0x4C$test_pe$test_opt_reg_a$__DOLLAR__procdff__DOLLAR__3625$reg0(.PORT_ID_ARST(fresh_wire_2224),
.PORT_ID_CLK(fresh_wire_2223),
.PORT_ID_IN(fresh_wire_2221),
.PORT_ID_OUT(fresh_wire_2222));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000011),
.PARAM_OUT_WIDTH(32'h00000022)) pe_0x4C$test_pe$test_pe_comp$test_mult_add$__DOLLAR__mul__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__1503$extendA(.PORT_ID_IN(fresh_wire_2225),
.PORT_ID_OUT(fresh_wire_2226));

	CELL_TYPE_MUL #(.PARAM_WIDTH(32'h00000022)) pe_0x4C$test_pe$test_pe_comp$test_mult_add$__DOLLAR__mul__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__1503$op0(.PORT_ID_IN0(fresh_wire_2227),
.PORT_ID_IN1(fresh_wire_2228),
.PORT_ID_OUT(fresh_wire_2229));

	CELL_TYPE_REG_ARST #(.PARAM_ARST_POSEDGE(1'h0),
.PARAM_CLK_POSEDGE(1'h1),
.PARAM_INIT_VALUE(16'h0000),
.PARAM_WIDTH(32'h00000010)) pe_0x57$test_pe$test_opt_reg_a$__DOLLAR__procdff__DOLLAR__3625$reg0(.PORT_ID_ARST(fresh_wire_2233),
.PORT_ID_CLK(fresh_wire_2232),
.PORT_ID_IN(fresh_wire_2230),
.PORT_ID_OUT(fresh_wire_2231));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000011),
.PARAM_OUT_WIDTH(32'h00000022)) pe_0x57$test_pe$test_pe_comp$test_mult_add$__DOLLAR__mul__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__1503$extendA(.PORT_ID_IN(fresh_wire_2234),
.PORT_ID_OUT(fresh_wire_2235));

	CELL_TYPE_MUL #(.PARAM_WIDTH(32'h00000022)) pe_0x57$test_pe$test_pe_comp$test_mult_add$__DOLLAR__mul__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__1503$op0(.PORT_ID_IN0(fresh_wire_2236),
.PORT_ID_IN1(fresh_wire_2237),
.PORT_ID_OUT(fresh_wire_2238));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000011)) pe_0x5A$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$extendA(.PORT_ID_IN(fresh_wire_2239),
.PORT_ID_OUT(fresh_wire_2240));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000010),
.PARAM_OUT_WIDTH(32'h00000011)) pe_0x5A$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$extendB(.PORT_ID_IN(fresh_wire_2241),
.PORT_ID_OUT(fresh_wire_2242));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000011)) pe_0x5A$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1494$op0(.PORT_ID_IN0(fresh_wire_2243),
.PORT_ID_IN1(fresh_wire_2244),
.PORT_ID_OUT(fresh_wire_2245));

	CELL_TYPE_ADD #(.PARAM_WIDTH(32'h00000011)) pe_0x5A$test_pe$test_pe_comp$GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add$__DOLLAR__add__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__1495$op0(.PORT_ID_IN0(fresh_wire_2246),
.PORT_ID_IN1(fresh_wire_2247),
.PORT_ID_OUT(fresh_wire_2248));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) pe_0xFF__DOT__tile_id__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(.PORT_ID_OUT(fresh_wire_2249));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) reset_in_port_cell(.PORT_ID_IN(reset_in),
.PORT_ID_OUT(fresh_wire_148));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) tck_port_cell(.PORT_ID_IN(tck),
.PORT_ID_OUT(fresh_wire_149));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) tdi_port_cell(.PORT_ID_IN(tdi),
.PORT_ID_OUT(fresh_wire_150));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) tdo_port_cell(.PORT_ID_IN(fresh_wire_151),
.PORT_ID_OUT(tdo));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) tms_port_cell(.PORT_ID_IN(tms),
.PORT_ID_OUT(fresh_wire_152));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) trst_n_port_cell(.PORT_ID_IN(trst_n),
.PORT_ID_OUT(fresh_wire_153));

	assign fresh_wire_0[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_13[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_14[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_15[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_16[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_17[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_18[ 0 ] = fresh_wire_154[ 0 ];
	assign fresh_wire_18[ 1 ] = fresh_wire_154[ 1 ];
	assign fresh_wire_18[ 2 ] = fresh_wire_154[ 2 ];
	assign fresh_wire_18[ 3 ] = fresh_wire_154[ 3 ];
	assign fresh_wire_18[ 4 ] = fresh_wire_154[ 4 ];
	assign fresh_wire_18[ 5 ] = fresh_wire_154[ 5 ];
	assign fresh_wire_18[ 6 ] = fresh_wire_154[ 6 ];
	assign fresh_wire_18[ 7 ] = fresh_wire_154[ 7 ];
	assign fresh_wire_18[ 8 ] = fresh_wire_154[ 8 ];
	assign fresh_wire_18[ 9 ] = fresh_wire_154[ 9 ];
	assign fresh_wire_18[ 10 ] = fresh_wire_154[ 10 ];
	assign fresh_wire_18[ 11 ] = fresh_wire_154[ 11 ];
	assign fresh_wire_18[ 12 ] = fresh_wire_154[ 12 ];
	assign fresh_wire_19[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_19[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_19[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_19[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_21[ 0 ] = fresh_wire_2215[ 15 ];
	assign fresh_wire_23[ 0 ] = fresh_wire_2215[ 5 ];
	assign fresh_wire_25[ 0 ] = fresh_wire_2215[ 4 ];
	assign fresh_wire_27[ 0 ] = fresh_wire_2215[ 3 ];
	assign fresh_wire_29[ 0 ] = fresh_wire_2215[ 2 ];
	assign fresh_wire_31[ 0 ] = fresh_wire_2215[ 1 ];
	assign fresh_wire_33[ 0 ] = fresh_wire_2215[ 0 ];
	assign fresh_wire_35[ 0 ] = fresh_wire_2215[ 14 ];
	assign fresh_wire_37[ 0 ] = fresh_wire_2215[ 13 ];
	assign fresh_wire_39[ 0 ] = fresh_wire_2215[ 12 ];
	assign fresh_wire_41[ 0 ] = fresh_wire_2215[ 11 ];
	assign fresh_wire_43[ 0 ] = fresh_wire_2215[ 10 ];
	assign fresh_wire_45[ 0 ] = fresh_wire_2215[ 9 ];
	assign fresh_wire_47[ 0 ] = fresh_wire_2215[ 8 ];
	assign fresh_wire_49[ 0 ] = fresh_wire_2215[ 7 ];
	assign fresh_wire_51[ 0 ] = fresh_wire_2215[ 6 ];
	assign fresh_wire_53[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_55[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_57[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_59[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_61[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_63[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_65[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_67[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_69[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_71[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_73[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_75[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_77[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_79[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_81[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_83[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_85[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_87[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_89[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_91[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_93[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_95[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_97[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_99[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_101[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_103[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_105[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_107[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_109[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_111[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_113[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_115[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_117[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_119[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_121[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_123[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_125[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_127[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_129[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_131[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_133[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_135[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_137[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_139[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_141[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_143[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_145[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_147[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_151[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_155[ 0 ] = fresh_wire_2117[ 0 ];
	assign fresh_wire_156[ 0 ] = fresh_wire_163[ 0 ];
	assign fresh_wire_158[ 0 ] = fresh_wire_2117[ 0 ];
	assign fresh_wire_159[ 0 ] = fresh_wire_163[ 0 ];
	assign fresh_wire_161[ 0 ] = fresh_wire_426[ 0 ];
	assign fresh_wire_162[ 0 ] = fresh_wire_201[ 0 ];
	assign fresh_wire_164[ 0 ] = fresh_wire_406[ 0 ];
	assign fresh_wire_164[ 1 ] = fresh_wire_406[ 1 ];
	assign fresh_wire_164[ 2 ] = fresh_wire_406[ 2 ];
	assign fresh_wire_164[ 3 ] = fresh_wire_406[ 3 ];
	assign fresh_wire_164[ 4 ] = fresh_wire_406[ 4 ];
	assign fresh_wire_164[ 5 ] = fresh_wire_406[ 5 ];
	assign fresh_wire_164[ 6 ] = fresh_wire_406[ 6 ];
	assign fresh_wire_164[ 7 ] = fresh_wire_406[ 7 ];
	assign fresh_wire_164[ 8 ] = fresh_wire_406[ 8 ];
	assign fresh_wire_164[ 9 ] = fresh_wire_406[ 9 ];
	assign fresh_wire_164[ 10 ] = fresh_wire_406[ 10 ];
	assign fresh_wire_164[ 11 ] = fresh_wire_406[ 11 ];
	assign fresh_wire_164[ 12 ] = fresh_wire_406[ 12 ];
	assign fresh_wire_164[ 13 ] = fresh_wire_406[ 13 ];
	assign fresh_wire_164[ 14 ] = fresh_wire_406[ 14 ];
	assign fresh_wire_164[ 15 ] = fresh_wire_406[ 15 ];
	assign fresh_wire_165[ 0 ] = fresh_wire_2251[ 0 ];
	assign fresh_wire_165[ 1 ] = fresh_wire_2251[ 1 ];
	assign fresh_wire_165[ 2 ] = fresh_wire_2251[ 2 ];
	assign fresh_wire_165[ 3 ] = fresh_wire_2251[ 3 ];
	assign fresh_wire_165[ 4 ] = fresh_wire_2251[ 4 ];
	assign fresh_wire_165[ 5 ] = fresh_wire_2251[ 5 ];
	assign fresh_wire_165[ 6 ] = fresh_wire_2251[ 6 ];
	assign fresh_wire_165[ 7 ] = fresh_wire_2251[ 7 ];
	assign fresh_wire_165[ 8 ] = fresh_wire_2251[ 8 ];
	assign fresh_wire_165[ 9 ] = fresh_wire_2251[ 9 ];
	assign fresh_wire_165[ 10 ] = fresh_wire_2251[ 10 ];
	assign fresh_wire_165[ 11 ] = fresh_wire_2251[ 11 ];
	assign fresh_wire_165[ 12 ] = fresh_wire_2251[ 12 ];
	assign fresh_wire_165[ 13 ] = fresh_wire_2251[ 13 ];
	assign fresh_wire_165[ 14 ] = fresh_wire_2251[ 14 ];
	assign fresh_wire_165[ 15 ] = fresh_wire_2251[ 15 ];
	assign fresh_wire_167[ 0 ] = fresh_wire_666[ 0 ];
	assign fresh_wire_167[ 1 ] = fresh_wire_666[ 1 ];
	assign fresh_wire_169[ 0 ] = fresh_wire_418[ 0 ];
	assign fresh_wire_169[ 1 ] = fresh_wire_418[ 1 ];
	assign fresh_wire_169[ 2 ] = fresh_wire_418[ 2 ];
	assign fresh_wire_169[ 3 ] = fresh_wire_418[ 3 ];
	assign fresh_wire_169[ 4 ] = fresh_wire_418[ 4 ];
	assign fresh_wire_169[ 5 ] = fresh_wire_418[ 5 ];
	assign fresh_wire_169[ 6 ] = fresh_wire_418[ 6 ];
	assign fresh_wire_169[ 7 ] = fresh_wire_418[ 7 ];
	assign fresh_wire_169[ 8 ] = fresh_wire_418[ 8 ];
	assign fresh_wire_169[ 9 ] = fresh_wire_418[ 9 ];
	assign fresh_wire_169[ 10 ] = fresh_wire_418[ 10 ];
	assign fresh_wire_169[ 11 ] = fresh_wire_418[ 11 ];
	assign fresh_wire_169[ 12 ] = fresh_wire_418[ 12 ];
	assign fresh_wire_169[ 13 ] = fresh_wire_418[ 13 ];
	assign fresh_wire_169[ 14 ] = fresh_wire_418[ 14 ];
	assign fresh_wire_169[ 15 ] = fresh_wire_418[ 15 ];
	assign fresh_wire_170[ 0 ] = fresh_wire_168[ 0 ];
	assign fresh_wire_170[ 1 ] = fresh_wire_168[ 1 ];
	assign fresh_wire_170[ 2 ] = fresh_wire_168[ 2 ];
	assign fresh_wire_170[ 3 ] = fresh_wire_168[ 3 ];
	assign fresh_wire_170[ 4 ] = fresh_wire_168[ 4 ];
	assign fresh_wire_170[ 5 ] = fresh_wire_168[ 5 ];
	assign fresh_wire_170[ 6 ] = fresh_wire_168[ 6 ];
	assign fresh_wire_170[ 7 ] = fresh_wire_168[ 7 ];
	assign fresh_wire_170[ 8 ] = fresh_wire_168[ 8 ];
	assign fresh_wire_170[ 9 ] = fresh_wire_168[ 9 ];
	assign fresh_wire_170[ 10 ] = fresh_wire_168[ 10 ];
	assign fresh_wire_170[ 11 ] = fresh_wire_168[ 11 ];
	assign fresh_wire_170[ 12 ] = fresh_wire_168[ 12 ];
	assign fresh_wire_170[ 13 ] = fresh_wire_168[ 13 ];
	assign fresh_wire_170[ 14 ] = fresh_wire_168[ 14 ];
	assign fresh_wire_170[ 15 ] = fresh_wire_168[ 15 ];
	assign fresh_wire_172[ 0 ] = fresh_wire_414[ 0 ];
	assign fresh_wire_172[ 1 ] = fresh_wire_414[ 1 ];
	assign fresh_wire_172[ 2 ] = fresh_wire_414[ 2 ];
	assign fresh_wire_172[ 3 ] = fresh_wire_414[ 3 ];
	assign fresh_wire_172[ 4 ] = fresh_wire_414[ 4 ];
	assign fresh_wire_172[ 5 ] = fresh_wire_414[ 5 ];
	assign fresh_wire_172[ 6 ] = fresh_wire_414[ 6 ];
	assign fresh_wire_172[ 7 ] = fresh_wire_414[ 7 ];
	assign fresh_wire_172[ 8 ] = fresh_wire_414[ 8 ];
	assign fresh_wire_172[ 9 ] = fresh_wire_414[ 9 ];
	assign fresh_wire_172[ 10 ] = fresh_wire_414[ 10 ];
	assign fresh_wire_172[ 11 ] = fresh_wire_414[ 11 ];
	assign fresh_wire_172[ 12 ] = fresh_wire_414[ 12 ];
	assign fresh_wire_172[ 13 ] = fresh_wire_414[ 13 ];
	assign fresh_wire_172[ 14 ] = fresh_wire_414[ 14 ];
	assign fresh_wire_172[ 15 ] = fresh_wire_414[ 15 ];
	assign fresh_wire_174[ 0 ] = fresh_wire_173[ 0 ];
	assign fresh_wire_174[ 1 ] = fresh_wire_173[ 1 ];
	assign fresh_wire_174[ 2 ] = fresh_wire_173[ 2 ];
	assign fresh_wire_174[ 3 ] = fresh_wire_173[ 3 ];
	assign fresh_wire_174[ 4 ] = fresh_wire_173[ 4 ];
	assign fresh_wire_174[ 5 ] = fresh_wire_173[ 5 ];
	assign fresh_wire_174[ 6 ] = fresh_wire_173[ 6 ];
	assign fresh_wire_174[ 7 ] = fresh_wire_173[ 7 ];
	assign fresh_wire_174[ 8 ] = fresh_wire_173[ 8 ];
	assign fresh_wire_174[ 9 ] = fresh_wire_173[ 9 ];
	assign fresh_wire_174[ 10 ] = fresh_wire_173[ 10 ];
	assign fresh_wire_174[ 11 ] = fresh_wire_173[ 11 ];
	assign fresh_wire_174[ 12 ] = fresh_wire_173[ 12 ];
	assign fresh_wire_174[ 13 ] = fresh_wire_173[ 13 ];
	assign fresh_wire_174[ 14 ] = fresh_wire_173[ 14 ];
	assign fresh_wire_174[ 15 ] = fresh_wire_173[ 15 ];
	assign fresh_wire_174[ 16 ] = fresh_wire_173[ 16 ];
	assign fresh_wire_174[ 17 ] = fresh_wire_173[ 17 ];
	assign fresh_wire_174[ 18 ] = fresh_wire_173[ 18 ];
	assign fresh_wire_174[ 19 ] = fresh_wire_173[ 19 ];
	assign fresh_wire_174[ 20 ] = fresh_wire_173[ 20 ];
	assign fresh_wire_174[ 21 ] = fresh_wire_173[ 21 ];
	assign fresh_wire_174[ 22 ] = fresh_wire_173[ 22 ];
	assign fresh_wire_174[ 23 ] = fresh_wire_173[ 23 ];
	assign fresh_wire_174[ 24 ] = fresh_wire_173[ 24 ];
	assign fresh_wire_174[ 25 ] = fresh_wire_173[ 25 ];
	assign fresh_wire_174[ 26 ] = fresh_wire_173[ 26 ];
	assign fresh_wire_174[ 27 ] = fresh_wire_173[ 27 ];
	assign fresh_wire_174[ 28 ] = fresh_wire_173[ 28 ];
	assign fresh_wire_174[ 29 ] = fresh_wire_173[ 29 ];
	assign fresh_wire_174[ 30 ] = fresh_wire_173[ 30 ];
	assign fresh_wire_174[ 31 ] = fresh_wire_173[ 31 ];
	assign fresh_wire_175[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_175[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 16 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 17 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 18 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 19 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 20 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 21 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 22 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 23 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 24 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 25 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 26 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 27 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 28 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 29 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 30 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_175[ 31 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_177[ 0 ] = fresh_wire_418[ 0 ];
	assign fresh_wire_177[ 1 ] = fresh_wire_418[ 1 ];
	assign fresh_wire_177[ 2 ] = fresh_wire_418[ 2 ];
	assign fresh_wire_177[ 3 ] = fresh_wire_418[ 3 ];
	assign fresh_wire_177[ 4 ] = fresh_wire_418[ 4 ];
	assign fresh_wire_177[ 5 ] = fresh_wire_418[ 5 ];
	assign fresh_wire_177[ 6 ] = fresh_wire_418[ 6 ];
	assign fresh_wire_177[ 7 ] = fresh_wire_418[ 7 ];
	assign fresh_wire_177[ 8 ] = fresh_wire_418[ 8 ];
	assign fresh_wire_177[ 9 ] = fresh_wire_418[ 9 ];
	assign fresh_wire_177[ 10 ] = fresh_wire_418[ 10 ];
	assign fresh_wire_177[ 11 ] = fresh_wire_418[ 11 ];
	assign fresh_wire_177[ 12 ] = fresh_wire_418[ 12 ];
	assign fresh_wire_177[ 13 ] = fresh_wire_418[ 13 ];
	assign fresh_wire_177[ 14 ] = fresh_wire_418[ 14 ];
	assign fresh_wire_177[ 15 ] = fresh_wire_418[ 15 ];
	assign fresh_wire_179[ 0 ] = fresh_wire_178[ 0 ];
	assign fresh_wire_179[ 1 ] = fresh_wire_178[ 1 ];
	assign fresh_wire_179[ 2 ] = fresh_wire_178[ 2 ];
	assign fresh_wire_179[ 3 ] = fresh_wire_178[ 3 ];
	assign fresh_wire_179[ 4 ] = fresh_wire_178[ 4 ];
	assign fresh_wire_179[ 5 ] = fresh_wire_178[ 5 ];
	assign fresh_wire_179[ 6 ] = fresh_wire_178[ 6 ];
	assign fresh_wire_179[ 7 ] = fresh_wire_178[ 7 ];
	assign fresh_wire_179[ 8 ] = fresh_wire_178[ 8 ];
	assign fresh_wire_179[ 9 ] = fresh_wire_178[ 9 ];
	assign fresh_wire_179[ 10 ] = fresh_wire_178[ 10 ];
	assign fresh_wire_179[ 11 ] = fresh_wire_178[ 11 ];
	assign fresh_wire_179[ 12 ] = fresh_wire_178[ 12 ];
	assign fresh_wire_179[ 13 ] = fresh_wire_178[ 13 ];
	assign fresh_wire_179[ 14 ] = fresh_wire_178[ 14 ];
	assign fresh_wire_179[ 15 ] = fresh_wire_178[ 15 ];
	assign fresh_wire_179[ 16 ] = fresh_wire_178[ 16 ];
	assign fresh_wire_179[ 17 ] = fresh_wire_178[ 17 ];
	assign fresh_wire_179[ 18 ] = fresh_wire_178[ 18 ];
	assign fresh_wire_179[ 19 ] = fresh_wire_178[ 19 ];
	assign fresh_wire_179[ 20 ] = fresh_wire_178[ 20 ];
	assign fresh_wire_179[ 21 ] = fresh_wire_178[ 21 ];
	assign fresh_wire_179[ 22 ] = fresh_wire_178[ 22 ];
	assign fresh_wire_179[ 23 ] = fresh_wire_178[ 23 ];
	assign fresh_wire_179[ 24 ] = fresh_wire_178[ 24 ];
	assign fresh_wire_179[ 25 ] = fresh_wire_178[ 25 ];
	assign fresh_wire_179[ 26 ] = fresh_wire_178[ 26 ];
	assign fresh_wire_179[ 27 ] = fresh_wire_178[ 27 ];
	assign fresh_wire_179[ 28 ] = fresh_wire_178[ 28 ];
	assign fresh_wire_179[ 29 ] = fresh_wire_178[ 29 ];
	assign fresh_wire_179[ 30 ] = fresh_wire_178[ 30 ];
	assign fresh_wire_179[ 31 ] = fresh_wire_178[ 31 ];
	assign fresh_wire_180[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 1 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_180[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 16 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 17 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 18 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 19 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 20 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 21 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 22 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 23 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 24 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 25 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 26 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 27 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 28 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 29 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 30 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_180[ 31 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_182[ 0 ] = fresh_wire_410[ 0 ];
	assign fresh_wire_182[ 1 ] = fresh_wire_410[ 1 ];
	assign fresh_wire_182[ 2 ] = fresh_wire_410[ 2 ];
	assign fresh_wire_182[ 3 ] = fresh_wire_410[ 3 ];
	assign fresh_wire_182[ 4 ] = fresh_wire_410[ 4 ];
	assign fresh_wire_182[ 5 ] = fresh_wire_410[ 5 ];
	assign fresh_wire_182[ 6 ] = fresh_wire_410[ 6 ];
	assign fresh_wire_182[ 7 ] = fresh_wire_410[ 7 ];
	assign fresh_wire_182[ 8 ] = fresh_wire_410[ 8 ];
	assign fresh_wire_182[ 9 ] = fresh_wire_410[ 9 ];
	assign fresh_wire_182[ 10 ] = fresh_wire_410[ 10 ];
	assign fresh_wire_182[ 11 ] = fresh_wire_410[ 11 ];
	assign fresh_wire_182[ 12 ] = fresh_wire_410[ 12 ];
	assign fresh_wire_182[ 13 ] = fresh_wire_410[ 13 ];
	assign fresh_wire_182[ 14 ] = fresh_wire_410[ 14 ];
	assign fresh_wire_182[ 15 ] = fresh_wire_410[ 15 ];
	assign fresh_wire_184[ 0 ] = fresh_wire_183[ 0 ];
	assign fresh_wire_184[ 1 ] = fresh_wire_183[ 1 ];
	assign fresh_wire_184[ 2 ] = fresh_wire_183[ 2 ];
	assign fresh_wire_184[ 3 ] = fresh_wire_183[ 3 ];
	assign fresh_wire_184[ 4 ] = fresh_wire_183[ 4 ];
	assign fresh_wire_184[ 5 ] = fresh_wire_183[ 5 ];
	assign fresh_wire_184[ 6 ] = fresh_wire_183[ 6 ];
	assign fresh_wire_184[ 7 ] = fresh_wire_183[ 7 ];
	assign fresh_wire_184[ 8 ] = fresh_wire_183[ 8 ];
	assign fresh_wire_184[ 9 ] = fresh_wire_183[ 9 ];
	assign fresh_wire_184[ 10 ] = fresh_wire_183[ 10 ];
	assign fresh_wire_184[ 11 ] = fresh_wire_183[ 11 ];
	assign fresh_wire_184[ 12 ] = fresh_wire_183[ 12 ];
	assign fresh_wire_184[ 13 ] = fresh_wire_183[ 13 ];
	assign fresh_wire_184[ 14 ] = fresh_wire_183[ 14 ];
	assign fresh_wire_184[ 15 ] = fresh_wire_183[ 15 ];
	assign fresh_wire_184[ 16 ] = fresh_wire_183[ 16 ];
	assign fresh_wire_184[ 17 ] = fresh_wire_183[ 17 ];
	assign fresh_wire_184[ 18 ] = fresh_wire_183[ 18 ];
	assign fresh_wire_184[ 19 ] = fresh_wire_183[ 19 ];
	assign fresh_wire_184[ 20 ] = fresh_wire_183[ 20 ];
	assign fresh_wire_184[ 21 ] = fresh_wire_183[ 21 ];
	assign fresh_wire_184[ 22 ] = fresh_wire_183[ 22 ];
	assign fresh_wire_184[ 23 ] = fresh_wire_183[ 23 ];
	assign fresh_wire_184[ 24 ] = fresh_wire_183[ 24 ];
	assign fresh_wire_184[ 25 ] = fresh_wire_183[ 25 ];
	assign fresh_wire_184[ 26 ] = fresh_wire_183[ 26 ];
	assign fresh_wire_184[ 27 ] = fresh_wire_183[ 27 ];
	assign fresh_wire_184[ 28 ] = fresh_wire_183[ 28 ];
	assign fresh_wire_184[ 29 ] = fresh_wire_183[ 29 ];
	assign fresh_wire_184[ 30 ] = fresh_wire_183[ 30 ];
	assign fresh_wire_184[ 31 ] = fresh_wire_183[ 31 ];
	assign fresh_wire_185[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_185[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 16 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 17 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 18 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 19 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 20 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 21 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 22 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 23 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 24 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 25 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 26 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 27 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 28 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 29 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 30 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_185[ 31 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_187[ 0 ] = fresh_wire_406[ 0 ];
	assign fresh_wire_187[ 1 ] = fresh_wire_406[ 1 ];
	assign fresh_wire_187[ 2 ] = fresh_wire_406[ 2 ];
	assign fresh_wire_187[ 3 ] = fresh_wire_406[ 3 ];
	assign fresh_wire_187[ 4 ] = fresh_wire_406[ 4 ];
	assign fresh_wire_187[ 5 ] = fresh_wire_406[ 5 ];
	assign fresh_wire_187[ 6 ] = fresh_wire_406[ 6 ];
	assign fresh_wire_187[ 7 ] = fresh_wire_406[ 7 ];
	assign fresh_wire_187[ 8 ] = fresh_wire_406[ 8 ];
	assign fresh_wire_187[ 9 ] = fresh_wire_406[ 9 ];
	assign fresh_wire_187[ 10 ] = fresh_wire_406[ 10 ];
	assign fresh_wire_187[ 11 ] = fresh_wire_406[ 11 ];
	assign fresh_wire_187[ 12 ] = fresh_wire_406[ 12 ];
	assign fresh_wire_187[ 13 ] = fresh_wire_406[ 13 ];
	assign fresh_wire_187[ 14 ] = fresh_wire_406[ 14 ];
	assign fresh_wire_187[ 15 ] = fresh_wire_406[ 15 ];
	assign fresh_wire_188[ 0 ] = fresh_wire_2252[ 0 ];
	assign fresh_wire_188[ 1 ] = fresh_wire_2252[ 1 ];
	assign fresh_wire_188[ 2 ] = fresh_wire_2252[ 2 ];
	assign fresh_wire_188[ 3 ] = fresh_wire_2252[ 3 ];
	assign fresh_wire_188[ 4 ] = fresh_wire_2252[ 4 ];
	assign fresh_wire_188[ 5 ] = fresh_wire_2252[ 5 ];
	assign fresh_wire_188[ 6 ] = fresh_wire_2252[ 6 ];
	assign fresh_wire_188[ 7 ] = fresh_wire_2252[ 7 ];
	assign fresh_wire_188[ 8 ] = fresh_wire_2252[ 8 ];
	assign fresh_wire_188[ 9 ] = fresh_wire_2252[ 9 ];
	assign fresh_wire_188[ 10 ] = fresh_wire_2252[ 10 ];
	assign fresh_wire_188[ 11 ] = fresh_wire_2252[ 11 ];
	assign fresh_wire_188[ 12 ] = fresh_wire_2252[ 12 ];
	assign fresh_wire_188[ 13 ] = fresh_wire_2252[ 13 ];
	assign fresh_wire_188[ 14 ] = fresh_wire_2252[ 14 ];
	assign fresh_wire_188[ 15 ] = fresh_wire_2252[ 15 ];
	assign fresh_wire_190[ 0 ] = fresh_wire_406[ 0 ];
	assign fresh_wire_190[ 1 ] = fresh_wire_406[ 1 ];
	assign fresh_wire_190[ 2 ] = fresh_wire_406[ 2 ];
	assign fresh_wire_190[ 3 ] = fresh_wire_406[ 3 ];
	assign fresh_wire_190[ 4 ] = fresh_wire_406[ 4 ];
	assign fresh_wire_190[ 5 ] = fresh_wire_406[ 5 ];
	assign fresh_wire_190[ 6 ] = fresh_wire_406[ 6 ];
	assign fresh_wire_190[ 7 ] = fresh_wire_406[ 7 ];
	assign fresh_wire_190[ 8 ] = fresh_wire_406[ 8 ];
	assign fresh_wire_190[ 9 ] = fresh_wire_406[ 9 ];
	assign fresh_wire_190[ 10 ] = fresh_wire_406[ 10 ];
	assign fresh_wire_190[ 11 ] = fresh_wire_406[ 11 ];
	assign fresh_wire_190[ 12 ] = fresh_wire_406[ 12 ];
	assign fresh_wire_190[ 13 ] = fresh_wire_406[ 13 ];
	assign fresh_wire_190[ 14 ] = fresh_wire_406[ 14 ];
	assign fresh_wire_190[ 15 ] = fresh_wire_406[ 15 ];
	assign fresh_wire_191[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_191[ 1 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_191[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_191[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_191[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_191[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_191[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_191[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_191[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_191[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_191[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_191[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_191[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_191[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_191[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_191[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_193[ 0 ] = fresh_wire_406[ 0 ];
	assign fresh_wire_193[ 1 ] = fresh_wire_406[ 1 ];
	assign fresh_wire_193[ 2 ] = fresh_wire_406[ 2 ];
	assign fresh_wire_193[ 3 ] = fresh_wire_406[ 3 ];
	assign fresh_wire_193[ 4 ] = fresh_wire_406[ 4 ];
	assign fresh_wire_193[ 5 ] = fresh_wire_406[ 5 ];
	assign fresh_wire_193[ 6 ] = fresh_wire_406[ 6 ];
	assign fresh_wire_193[ 7 ] = fresh_wire_406[ 7 ];
	assign fresh_wire_193[ 8 ] = fresh_wire_406[ 8 ];
	assign fresh_wire_193[ 9 ] = fresh_wire_406[ 9 ];
	assign fresh_wire_193[ 10 ] = fresh_wire_406[ 10 ];
	assign fresh_wire_193[ 11 ] = fresh_wire_406[ 11 ];
	assign fresh_wire_193[ 12 ] = fresh_wire_406[ 12 ];
	assign fresh_wire_193[ 13 ] = fresh_wire_406[ 13 ];
	assign fresh_wire_193[ 14 ] = fresh_wire_406[ 14 ];
	assign fresh_wire_193[ 15 ] = fresh_wire_406[ 15 ];
	assign fresh_wire_194[ 0 ] = fresh_wire_2253[ 0 ];
	assign fresh_wire_194[ 1 ] = fresh_wire_2253[ 1 ];
	assign fresh_wire_194[ 2 ] = fresh_wire_2253[ 2 ];
	assign fresh_wire_194[ 3 ] = fresh_wire_2253[ 3 ];
	assign fresh_wire_194[ 4 ] = fresh_wire_2253[ 4 ];
	assign fresh_wire_194[ 5 ] = fresh_wire_2253[ 5 ];
	assign fresh_wire_194[ 6 ] = fresh_wire_2253[ 6 ];
	assign fresh_wire_194[ 7 ] = fresh_wire_2253[ 7 ];
	assign fresh_wire_194[ 8 ] = fresh_wire_2253[ 8 ];
	assign fresh_wire_194[ 9 ] = fresh_wire_2253[ 9 ];
	assign fresh_wire_194[ 10 ] = fresh_wire_2253[ 10 ];
	assign fresh_wire_194[ 11 ] = fresh_wire_2253[ 11 ];
	assign fresh_wire_194[ 12 ] = fresh_wire_2253[ 12 ];
	assign fresh_wire_194[ 13 ] = fresh_wire_2253[ 13 ];
	assign fresh_wire_194[ 14 ] = fresh_wire_2253[ 14 ];
	assign fresh_wire_194[ 15 ] = fresh_wire_2253[ 15 ];
	assign fresh_wire_196[ 0 ] = fresh_wire_406[ 0 ];
	assign fresh_wire_196[ 1 ] = fresh_wire_406[ 1 ];
	assign fresh_wire_196[ 2 ] = fresh_wire_406[ 2 ];
	assign fresh_wire_196[ 3 ] = fresh_wire_406[ 3 ];
	assign fresh_wire_196[ 4 ] = fresh_wire_406[ 4 ];
	assign fresh_wire_196[ 5 ] = fresh_wire_406[ 5 ];
	assign fresh_wire_196[ 6 ] = fresh_wire_406[ 6 ];
	assign fresh_wire_196[ 7 ] = fresh_wire_406[ 7 ];
	assign fresh_wire_196[ 8 ] = fresh_wire_406[ 8 ];
	assign fresh_wire_196[ 9 ] = fresh_wire_406[ 9 ];
	assign fresh_wire_196[ 10 ] = fresh_wire_406[ 10 ];
	assign fresh_wire_196[ 11 ] = fresh_wire_406[ 11 ];
	assign fresh_wire_196[ 12 ] = fresh_wire_406[ 12 ];
	assign fresh_wire_196[ 13 ] = fresh_wire_406[ 13 ];
	assign fresh_wire_196[ 14 ] = fresh_wire_406[ 14 ];
	assign fresh_wire_196[ 15 ] = fresh_wire_406[ 15 ];
	assign fresh_wire_197[ 0 ] = fresh_wire_2254[ 0 ];
	assign fresh_wire_197[ 1 ] = fresh_wire_2254[ 1 ];
	assign fresh_wire_197[ 2 ] = fresh_wire_2254[ 2 ];
	assign fresh_wire_197[ 3 ] = fresh_wire_2254[ 3 ];
	assign fresh_wire_197[ 4 ] = fresh_wire_2254[ 4 ];
	assign fresh_wire_197[ 5 ] = fresh_wire_2254[ 5 ];
	assign fresh_wire_197[ 6 ] = fresh_wire_2254[ 6 ];
	assign fresh_wire_197[ 7 ] = fresh_wire_2254[ 7 ];
	assign fresh_wire_197[ 8 ] = fresh_wire_2254[ 8 ];
	assign fresh_wire_197[ 9 ] = fresh_wire_2254[ 9 ];
	assign fresh_wire_197[ 10 ] = fresh_wire_2254[ 10 ];
	assign fresh_wire_197[ 11 ] = fresh_wire_2254[ 11 ];
	assign fresh_wire_197[ 12 ] = fresh_wire_2254[ 12 ];
	assign fresh_wire_197[ 13 ] = fresh_wire_2254[ 13 ];
	assign fresh_wire_197[ 14 ] = fresh_wire_2254[ 14 ];
	assign fresh_wire_197[ 15 ] = fresh_wire_2254[ 15 ];
	assign fresh_wire_199[ 0 ] = fresh_wire_219[ 0 ];
	assign fresh_wire_200[ 0 ] = fresh_wire_228[ 0 ];
	assign fresh_wire_202[ 0 ] = fresh_wire_376[ 0 ];
	assign fresh_wire_202[ 1 ] = fresh_wire_376[ 1 ];
	assign fresh_wire_203[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_203[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_205[ 0 ] = fresh_wire_373[ 0 ];
	assign fresh_wire_205[ 1 ] = fresh_wire_373[ 1 ];
	assign fresh_wire_206[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_206[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_208[ 0 ] = fresh_wire_666[ 0 ];
	assign fresh_wire_208[ 1 ] = fresh_wire_666[ 1 ];
	assign fresh_wire_209[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_209[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_211[ 0 ] = fresh_wire_166[ 0 ];
	assign fresh_wire_211[ 1 ] = fresh_wire_166[ 1 ];
	assign fresh_wire_211[ 2 ] = fresh_wire_166[ 2 ];
	assign fresh_wire_211[ 3 ] = fresh_wire_166[ 3 ];
	assign fresh_wire_211[ 4 ] = fresh_wire_166[ 4 ];
	assign fresh_wire_211[ 5 ] = fresh_wire_166[ 5 ];
	assign fresh_wire_211[ 6 ] = fresh_wire_166[ 6 ];
	assign fresh_wire_211[ 7 ] = fresh_wire_166[ 7 ];
	assign fresh_wire_211[ 8 ] = fresh_wire_166[ 8 ];
	assign fresh_wire_211[ 9 ] = fresh_wire_166[ 9 ];
	assign fresh_wire_211[ 10 ] = fresh_wire_166[ 10 ];
	assign fresh_wire_211[ 11 ] = fresh_wire_166[ 11 ];
	assign fresh_wire_211[ 12 ] = fresh_wire_166[ 12 ];
	assign fresh_wire_211[ 13 ] = fresh_wire_166[ 13 ];
	assign fresh_wire_211[ 14 ] = fresh_wire_166[ 14 ];
	assign fresh_wire_211[ 15 ] = fresh_wire_166[ 15 ];
	assign fresh_wire_212[ 0 ] = fresh_wire_2255[ 0 ];
	assign fresh_wire_212[ 1 ] = fresh_wire_2255[ 1 ];
	assign fresh_wire_212[ 2 ] = fresh_wire_2255[ 2 ];
	assign fresh_wire_212[ 3 ] = fresh_wire_2255[ 3 ];
	assign fresh_wire_212[ 4 ] = fresh_wire_2255[ 4 ];
	assign fresh_wire_212[ 5 ] = fresh_wire_2255[ 5 ];
	assign fresh_wire_212[ 6 ] = fresh_wire_2255[ 6 ];
	assign fresh_wire_212[ 7 ] = fresh_wire_2255[ 7 ];
	assign fresh_wire_212[ 8 ] = fresh_wire_2255[ 8 ];
	assign fresh_wire_212[ 9 ] = fresh_wire_2255[ 9 ];
	assign fresh_wire_212[ 10 ] = fresh_wire_2255[ 10 ];
	assign fresh_wire_212[ 11 ] = fresh_wire_2255[ 11 ];
	assign fresh_wire_212[ 12 ] = fresh_wire_2255[ 12 ];
	assign fresh_wire_212[ 13 ] = fresh_wire_2255[ 13 ];
	assign fresh_wire_212[ 14 ] = fresh_wire_2255[ 14 ];
	assign fresh_wire_212[ 15 ] = fresh_wire_2255[ 15 ];
	assign fresh_wire_214[ 0 ] = fresh_wire_422[ 0 ];
	assign fresh_wire_215[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_217[ 0 ] = fresh_wire_430[ 0 ];
	assign fresh_wire_218[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_220[ 0 ] = fresh_wire_678[ 0 ];
	assign fresh_wire_221[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_223[ 0 ] = fresh_wire_286[ 0 ];
	assign fresh_wire_224[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_226[ 0 ] = fresh_wire_402[ 0 ];
	assign fresh_wire_226[ 1 ] = fresh_wire_402[ 1 ];
	assign fresh_wire_227[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_227[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_229[ 0 ] = fresh_wire_430[ 0 ];
	assign fresh_wire_230[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_232[ 0 ] = fresh_wire_426[ 0 ];
	assign fresh_wire_233[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_235[ 0 ] = fresh_wire_402[ 0 ];
	assign fresh_wire_235[ 1 ] = fresh_wire_402[ 1 ];
	assign fresh_wire_236[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_236[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_238[ 0 ] = fresh_wire_363[ 0 ];
	assign fresh_wire_239[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_241[ 0 ] = fresh_wire_398[ 0 ];
	assign fresh_wire_242[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_244[ 0 ] = fresh_wire_402[ 0 ];
	assign fresh_wire_244[ 1 ] = fresh_wire_402[ 1 ];
	assign fresh_wire_245[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_245[ 1 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_247[ 0 ] = fresh_wire_373[ 0 ];
	assign fresh_wire_247[ 1 ] = fresh_wire_373[ 1 ];
	assign fresh_wire_248[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_248[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_250[ 0 ] = fresh_wire_198[ 0 ];
	assign fresh_wire_250[ 1 ] = fresh_wire_198[ 1 ];
	assign fresh_wire_250[ 2 ] = fresh_wire_198[ 2 ];
	assign fresh_wire_250[ 3 ] = fresh_wire_198[ 3 ];
	assign fresh_wire_250[ 4 ] = fresh_wire_198[ 4 ];
	assign fresh_wire_250[ 5 ] = fresh_wire_198[ 5 ];
	assign fresh_wire_250[ 6 ] = fresh_wire_198[ 6 ];
	assign fresh_wire_250[ 7 ] = fresh_wire_198[ 7 ];
	assign fresh_wire_250[ 8 ] = fresh_wire_198[ 8 ];
	assign fresh_wire_250[ 9 ] = fresh_wire_198[ 9 ];
	assign fresh_wire_250[ 10 ] = fresh_wire_198[ 10 ];
	assign fresh_wire_250[ 11 ] = fresh_wire_198[ 11 ];
	assign fresh_wire_250[ 12 ] = fresh_wire_198[ 12 ];
	assign fresh_wire_250[ 13 ] = fresh_wire_198[ 13 ];
	assign fresh_wire_250[ 14 ] = fresh_wire_198[ 14 ];
	assign fresh_wire_250[ 15 ] = fresh_wire_198[ 15 ];
	assign fresh_wire_251[ 0 ] = fresh_wire_2256[ 0 ];
	assign fresh_wire_251[ 1 ] = fresh_wire_2256[ 1 ];
	assign fresh_wire_251[ 2 ] = fresh_wire_2256[ 2 ];
	assign fresh_wire_251[ 3 ] = fresh_wire_2256[ 3 ];
	assign fresh_wire_251[ 4 ] = fresh_wire_2256[ 4 ];
	assign fresh_wire_251[ 5 ] = fresh_wire_2256[ 5 ];
	assign fresh_wire_251[ 6 ] = fresh_wire_2256[ 6 ];
	assign fresh_wire_251[ 7 ] = fresh_wire_2256[ 7 ];
	assign fresh_wire_251[ 8 ] = fresh_wire_2256[ 8 ];
	assign fresh_wire_251[ 9 ] = fresh_wire_2256[ 9 ];
	assign fresh_wire_251[ 10 ] = fresh_wire_2256[ 10 ];
	assign fresh_wire_251[ 11 ] = fresh_wire_2256[ 11 ];
	assign fresh_wire_251[ 12 ] = fresh_wire_2256[ 12 ];
	assign fresh_wire_251[ 13 ] = fresh_wire_2256[ 13 ];
	assign fresh_wire_251[ 14 ] = fresh_wire_2256[ 14 ];
	assign fresh_wire_251[ 15 ] = fresh_wire_2256[ 15 ];
	assign fresh_wire_253[ 0 ] = fresh_wire_894[ 0 ];
	assign fresh_wire_254[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_256[ 0 ] = fresh_wire_394[ 0 ];
	assign fresh_wire_257[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_259[ 0 ] = fresh_wire_414[ 0 ];
	assign fresh_wire_259[ 1 ] = fresh_wire_414[ 1 ];
	assign fresh_wire_259[ 2 ] = fresh_wire_414[ 2 ];
	assign fresh_wire_259[ 3 ] = fresh_wire_414[ 3 ];
	assign fresh_wire_259[ 4 ] = fresh_wire_414[ 4 ];
	assign fresh_wire_259[ 5 ] = fresh_wire_414[ 5 ];
	assign fresh_wire_259[ 6 ] = fresh_wire_414[ 6 ];
	assign fresh_wire_259[ 7 ] = fresh_wire_414[ 7 ];
	assign fresh_wire_259[ 8 ] = fresh_wire_414[ 8 ];
	assign fresh_wire_259[ 9 ] = fresh_wire_414[ 9 ];
	assign fresh_wire_259[ 10 ] = fresh_wire_414[ 10 ];
	assign fresh_wire_259[ 11 ] = fresh_wire_414[ 11 ];
	assign fresh_wire_259[ 12 ] = fresh_wire_414[ 12 ];
	assign fresh_wire_259[ 13 ] = fresh_wire_414[ 13 ];
	assign fresh_wire_259[ 14 ] = fresh_wire_414[ 14 ];
	assign fresh_wire_259[ 15 ] = fresh_wire_414[ 15 ];
	assign fresh_wire_260[ 0 ] = fresh_wire_2258[ 0 ];
	assign fresh_wire_260[ 1 ] = fresh_wire_2258[ 1 ];
	assign fresh_wire_260[ 2 ] = fresh_wire_2258[ 2 ];
	assign fresh_wire_260[ 3 ] = fresh_wire_2258[ 3 ];
	assign fresh_wire_260[ 4 ] = fresh_wire_2258[ 4 ];
	assign fresh_wire_260[ 5 ] = fresh_wire_2258[ 5 ];
	assign fresh_wire_260[ 6 ] = fresh_wire_2258[ 6 ];
	assign fresh_wire_260[ 7 ] = fresh_wire_2258[ 7 ];
	assign fresh_wire_260[ 8 ] = fresh_wire_2258[ 8 ];
	assign fresh_wire_260[ 9 ] = fresh_wire_2258[ 9 ];
	assign fresh_wire_260[ 10 ] = fresh_wire_2258[ 10 ];
	assign fresh_wire_260[ 11 ] = fresh_wire_2258[ 11 ];
	assign fresh_wire_260[ 12 ] = fresh_wire_2258[ 12 ];
	assign fresh_wire_260[ 13 ] = fresh_wire_2258[ 13 ];
	assign fresh_wire_260[ 14 ] = fresh_wire_2258[ 14 ];
	assign fresh_wire_260[ 15 ] = fresh_wire_2258[ 15 ];
	assign fresh_wire_262[ 0 ] = fresh_wire_410[ 0 ];
	assign fresh_wire_262[ 1 ] = fresh_wire_410[ 1 ];
	assign fresh_wire_262[ 2 ] = fresh_wire_410[ 2 ];
	assign fresh_wire_262[ 3 ] = fresh_wire_410[ 3 ];
	assign fresh_wire_262[ 4 ] = fresh_wire_410[ 4 ];
	assign fresh_wire_262[ 5 ] = fresh_wire_410[ 5 ];
	assign fresh_wire_262[ 6 ] = fresh_wire_410[ 6 ];
	assign fresh_wire_262[ 7 ] = fresh_wire_410[ 7 ];
	assign fresh_wire_262[ 8 ] = fresh_wire_410[ 8 ];
	assign fresh_wire_262[ 9 ] = fresh_wire_410[ 9 ];
	assign fresh_wire_262[ 10 ] = fresh_wire_410[ 10 ];
	assign fresh_wire_262[ 11 ] = fresh_wire_410[ 11 ];
	assign fresh_wire_262[ 12 ] = fresh_wire_410[ 12 ];
	assign fresh_wire_262[ 13 ] = fresh_wire_410[ 13 ];
	assign fresh_wire_262[ 14 ] = fresh_wire_410[ 14 ];
	assign fresh_wire_262[ 15 ] = fresh_wire_410[ 15 ];
	assign fresh_wire_263[ 0 ] = fresh_wire_2258[ 0 ];
	assign fresh_wire_263[ 1 ] = fresh_wire_2258[ 1 ];
	assign fresh_wire_263[ 2 ] = fresh_wire_2258[ 2 ];
	assign fresh_wire_263[ 3 ] = fresh_wire_2258[ 3 ];
	assign fresh_wire_263[ 4 ] = fresh_wire_2258[ 4 ];
	assign fresh_wire_263[ 5 ] = fresh_wire_2258[ 5 ];
	assign fresh_wire_263[ 6 ] = fresh_wire_2258[ 6 ];
	assign fresh_wire_263[ 7 ] = fresh_wire_2258[ 7 ];
	assign fresh_wire_263[ 8 ] = fresh_wire_2258[ 8 ];
	assign fresh_wire_263[ 9 ] = fresh_wire_2258[ 9 ];
	assign fresh_wire_263[ 10 ] = fresh_wire_2258[ 10 ];
	assign fresh_wire_263[ 11 ] = fresh_wire_2258[ 11 ];
	assign fresh_wire_263[ 12 ] = fresh_wire_2258[ 12 ];
	assign fresh_wire_263[ 13 ] = fresh_wire_2258[ 13 ];
	assign fresh_wire_263[ 14 ] = fresh_wire_2258[ 14 ];
	assign fresh_wire_263[ 15 ] = fresh_wire_2258[ 15 ];
	assign fresh_wire_265[ 0 ] = fresh_wire_195[ 0 ];
	assign fresh_wire_265[ 1 ] = fresh_wire_195[ 1 ];
	assign fresh_wire_265[ 2 ] = fresh_wire_195[ 2 ];
	assign fresh_wire_265[ 3 ] = fresh_wire_195[ 3 ];
	assign fresh_wire_265[ 4 ] = fresh_wire_195[ 4 ];
	assign fresh_wire_265[ 5 ] = fresh_wire_195[ 5 ];
	assign fresh_wire_265[ 6 ] = fresh_wire_195[ 6 ];
	assign fresh_wire_265[ 7 ] = fresh_wire_195[ 7 ];
	assign fresh_wire_265[ 8 ] = fresh_wire_195[ 8 ];
	assign fresh_wire_265[ 9 ] = fresh_wire_195[ 9 ];
	assign fresh_wire_265[ 10 ] = fresh_wire_195[ 10 ];
	assign fresh_wire_265[ 11 ] = fresh_wire_195[ 11 ];
	assign fresh_wire_265[ 12 ] = fresh_wire_195[ 12 ];
	assign fresh_wire_265[ 13 ] = fresh_wire_195[ 13 ];
	assign fresh_wire_265[ 14 ] = fresh_wire_195[ 14 ];
	assign fresh_wire_265[ 15 ] = fresh_wire_195[ 15 ];
	assign fresh_wire_266[ 0 ] = fresh_wire_2257[ 0 ];
	assign fresh_wire_266[ 1 ] = fresh_wire_2257[ 1 ];
	assign fresh_wire_266[ 2 ] = fresh_wire_2257[ 2 ];
	assign fresh_wire_266[ 3 ] = fresh_wire_2257[ 3 ];
	assign fresh_wire_266[ 4 ] = fresh_wire_2257[ 4 ];
	assign fresh_wire_266[ 5 ] = fresh_wire_2257[ 5 ];
	assign fresh_wire_266[ 6 ] = fresh_wire_2257[ 6 ];
	assign fresh_wire_266[ 7 ] = fresh_wire_2257[ 7 ];
	assign fresh_wire_266[ 8 ] = fresh_wire_2257[ 8 ];
	assign fresh_wire_266[ 9 ] = fresh_wire_2257[ 9 ];
	assign fresh_wire_266[ 10 ] = fresh_wire_2257[ 10 ];
	assign fresh_wire_266[ 11 ] = fresh_wire_2257[ 11 ];
	assign fresh_wire_266[ 12 ] = fresh_wire_2257[ 12 ];
	assign fresh_wire_266[ 13 ] = fresh_wire_2257[ 13 ];
	assign fresh_wire_266[ 14 ] = fresh_wire_2257[ 14 ];
	assign fresh_wire_266[ 15 ] = fresh_wire_2257[ 15 ];
	assign fresh_wire_268[ 0 ] = fresh_wire_204[ 0 ];
	assign fresh_wire_270[ 0 ] = fresh_wire_269[ 0 ];
	assign fresh_wire_271[ 0 ] = fresh_wire_274[ 0 ];
	assign fresh_wire_273[ 0 ] = fresh_wire_207[ 0 ];
	assign fresh_wire_275[ 0 ] = fresh_wire_272[ 0 ];
	assign fresh_wire_277[ 0 ] = fresh_wire_276[ 0 ];
	assign fresh_wire_278[ 0 ] = fresh_wire_281[ 0 ];
	assign fresh_wire_280[ 0 ] = fresh_wire_210[ 0 ];
	assign fresh_wire_282[ 0 ] = fresh_wire_279[ 0 ];
	assign fresh_wire_284[ 0 ] = fresh_wire_283[ 0 ];
	assign fresh_wire_285[ 0 ] = fresh_wire_288[ 0 ];
	assign fresh_wire_287[ 0 ] = fresh_wire_213[ 0 ];
	assign fresh_wire_289[ 0 ] = fresh_wire_237[ 0 ];
	assign fresh_wire_291[ 0 ] = fresh_wire_290[ 0 ];
	assign fresh_wire_292[ 0 ] = fresh_wire_2308[ 0 ];
	assign fresh_wire_294[ 0 ] = fresh_wire_293[ 0 ];
	assign fresh_wire_296[ 0 ] = fresh_wire_295[ 0 ];
	assign fresh_wire_297[ 0 ] = fresh_wire_300[ 0 ];
	assign fresh_wire_299[ 0 ] = fresh_wire_240[ 0 ];
	assign fresh_wire_301[ 0 ] = fresh_wire_228[ 0 ];
	assign fresh_wire_303[ 0 ] = fresh_wire_302[ 0 ];
	assign fresh_wire_304[ 0 ] = fresh_wire_2309[ 0 ];
	assign fresh_wire_306[ 0 ] = fresh_wire_305[ 0 ];
	assign fresh_wire_308[ 0 ] = fresh_wire_307[ 0 ];
	assign fresh_wire_309[ 0 ] = fresh_wire_312[ 0 ];
	assign fresh_wire_311[ 0 ] = fresh_wire_366[ 0 ];
	assign fresh_wire_313[ 0 ] = fresh_wire_228[ 0 ];
	assign fresh_wire_315[ 0 ] = fresh_wire_314[ 0 ];
	assign fresh_wire_316[ 0 ] = fresh_wire_319[ 0 ];
	assign fresh_wire_318[ 0 ] = fresh_wire_267[ 0 ];
	assign fresh_wire_320[ 0 ] = fresh_wire_2310[ 0 ];
	assign fresh_wire_321[ 0 ] = fresh_wire_324[ 0 ];
	assign fresh_wire_323[ 0 ] = fresh_wire_240[ 0 ];
	assign fresh_wire_325[ 0 ] = fresh_wire_246[ 0 ];
	assign fresh_wire_327[ 0 ] = fresh_wire_326[ 0 ];
	assign fresh_wire_328[ 0 ] = fresh_wire_2311[ 0 ];
	assign fresh_wire_330[ 0 ] = fresh_wire_204[ 0 ];
	assign fresh_wire_332[ 0 ] = fresh_wire_331[ 0 ];
	assign fresh_wire_333[ 0 ] = fresh_wire_336[ 0 ];
	assign fresh_wire_335[ 0 ] = fresh_wire_207[ 0 ];
	assign fresh_wire_337[ 0 ] = fresh_wire_334[ 0 ];
	assign fresh_wire_339[ 0 ] = fresh_wire_338[ 0 ];
	assign fresh_wire_340[ 0 ] = fresh_wire_343[ 0 ];
	assign fresh_wire_342[ 0 ] = fresh_wire_210[ 0 ];
	assign fresh_wire_344[ 0 ] = fresh_wire_341[ 0 ];
	assign fresh_wire_346[ 0 ] = fresh_wire_345[ 0 ];
	assign fresh_wire_347[ 0 ] = fresh_wire_350[ 0 ];
	assign fresh_wire_349[ 0 ] = fresh_wire_252[ 0 ];
	assign fresh_wire_351[ 0 ] = fresh_wire_255[ 0 ];
	assign fresh_wire_353[ 0 ] = fresh_wire_352[ 0 ];
	assign fresh_wire_354[ 0 ] = fresh_wire_2312[ 0 ];
	assign fresh_wire_356[ 0 ] = fresh_wire_363[ 0 ];
	assign fresh_wire_358[ 0 ] = fresh_wire_2313[ 0 ];
	assign fresh_wire_359[ 0 ] = fresh_wire_357[ 0 ];
	assign fresh_wire_361[ 0 ] = fresh_wire_171[ 0 ];
	assign fresh_wire_361[ 1 ] = fresh_wire_171[ 1 ];
	assign fresh_wire_361[ 2 ] = fresh_wire_171[ 2 ];
	assign fresh_wire_361[ 3 ] = fresh_wire_171[ 3 ];
	assign fresh_wire_361[ 4 ] = fresh_wire_171[ 4 ];
	assign fresh_wire_361[ 5 ] = fresh_wire_171[ 5 ];
	assign fresh_wire_361[ 6 ] = fresh_wire_171[ 6 ];
	assign fresh_wire_361[ 7 ] = fresh_wire_171[ 7 ];
	assign fresh_wire_361[ 8 ] = fresh_wire_171[ 8 ];
	assign fresh_wire_361[ 9 ] = fresh_wire_171[ 9 ];
	assign fresh_wire_361[ 10 ] = fresh_wire_171[ 10 ];
	assign fresh_wire_361[ 11 ] = fresh_wire_171[ 11 ];
	assign fresh_wire_361[ 12 ] = fresh_wire_171[ 12 ];
	assign fresh_wire_361[ 13 ] = fresh_wire_171[ 13 ];
	assign fresh_wire_361[ 14 ] = fresh_wire_171[ 14 ];
	assign fresh_wire_361[ 15 ] = fresh_wire_171[ 15 ];
	assign fresh_wire_362[ 0 ] = fresh_wire_2259[ 0 ];
	assign fresh_wire_362[ 1 ] = fresh_wire_2259[ 1 ];
	assign fresh_wire_362[ 2 ] = fresh_wire_2259[ 2 ];
	assign fresh_wire_362[ 3 ] = fresh_wire_2259[ 3 ];
	assign fresh_wire_362[ 4 ] = fresh_wire_2259[ 4 ];
	assign fresh_wire_362[ 5 ] = fresh_wire_2259[ 5 ];
	assign fresh_wire_362[ 6 ] = fresh_wire_2259[ 6 ];
	assign fresh_wire_362[ 7 ] = fresh_wire_2259[ 7 ];
	assign fresh_wire_362[ 8 ] = fresh_wire_2259[ 8 ];
	assign fresh_wire_362[ 9 ] = fresh_wire_2259[ 9 ];
	assign fresh_wire_362[ 10 ] = fresh_wire_2259[ 10 ];
	assign fresh_wire_362[ 11 ] = fresh_wire_2259[ 11 ];
	assign fresh_wire_362[ 12 ] = fresh_wire_2259[ 12 ];
	assign fresh_wire_362[ 13 ] = fresh_wire_2259[ 13 ];
	assign fresh_wire_362[ 14 ] = fresh_wire_2259[ 14 ];
	assign fresh_wire_362[ 15 ] = fresh_wire_2259[ 15 ];
	assign fresh_wire_364[ 0 ] = fresh_wire_189[ 0 ];
	assign fresh_wire_364[ 1 ] = fresh_wire_189[ 1 ];
	assign fresh_wire_364[ 2 ] = fresh_wire_189[ 2 ];
	assign fresh_wire_364[ 3 ] = fresh_wire_189[ 3 ];
	assign fresh_wire_364[ 4 ] = fresh_wire_189[ 4 ];
	assign fresh_wire_364[ 5 ] = fresh_wire_189[ 5 ];
	assign fresh_wire_364[ 6 ] = fresh_wire_189[ 6 ];
	assign fresh_wire_364[ 7 ] = fresh_wire_189[ 7 ];
	assign fresh_wire_364[ 8 ] = fresh_wire_189[ 8 ];
	assign fresh_wire_364[ 9 ] = fresh_wire_189[ 9 ];
	assign fresh_wire_364[ 10 ] = fresh_wire_189[ 10 ];
	assign fresh_wire_364[ 11 ] = fresh_wire_189[ 11 ];
	assign fresh_wire_364[ 12 ] = fresh_wire_189[ 12 ];
	assign fresh_wire_364[ 13 ] = fresh_wire_189[ 13 ];
	assign fresh_wire_364[ 14 ] = fresh_wire_189[ 14 ];
	assign fresh_wire_364[ 15 ] = fresh_wire_189[ 15 ];
	assign fresh_wire_365[ 0 ] = fresh_wire_2257[ 0 ];
	assign fresh_wire_365[ 1 ] = fresh_wire_2257[ 1 ];
	assign fresh_wire_365[ 2 ] = fresh_wire_2257[ 2 ];
	assign fresh_wire_365[ 3 ] = fresh_wire_2257[ 3 ];
	assign fresh_wire_365[ 4 ] = fresh_wire_2257[ 4 ];
	assign fresh_wire_365[ 5 ] = fresh_wire_2257[ 5 ];
	assign fresh_wire_365[ 6 ] = fresh_wire_2257[ 6 ];
	assign fresh_wire_365[ 7 ] = fresh_wire_2257[ 7 ];
	assign fresh_wire_365[ 8 ] = fresh_wire_2257[ 8 ];
	assign fresh_wire_365[ 9 ] = fresh_wire_2257[ 9 ];
	assign fresh_wire_365[ 10 ] = fresh_wire_2257[ 10 ];
	assign fresh_wire_365[ 11 ] = fresh_wire_2257[ 11 ];
	assign fresh_wire_365[ 12 ] = fresh_wire_2257[ 12 ];
	assign fresh_wire_365[ 13 ] = fresh_wire_2257[ 13 ];
	assign fresh_wire_365[ 14 ] = fresh_wire_2257[ 14 ];
	assign fresh_wire_365[ 15 ] = fresh_wire_2257[ 15 ];
	assign fresh_wire_367[ 0 ] = fresh_wire_430[ 0 ];
	assign fresh_wire_369[ 0 ] = fresh_wire_360[ 0 ];
	assign fresh_wire_371[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_372[ 0 ] = fresh_wire_402[ 0 ];
	assign fresh_wire_372[ 1 ] = fresh_wire_402[ 1 ];
	assign fresh_wire_374[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_375[ 0 ] = fresh_wire_373[ 0 ];
	assign fresh_wire_375[ 1 ] = fresh_wire_373[ 1 ];
	assign fresh_wire_377[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_378[ 0 ] = fresh_wire_878[ 0 ];
	assign fresh_wire_378[ 1 ] = fresh_wire_878[ 1 ];
	assign fresh_wire_378[ 2 ] = fresh_wire_878[ 2 ];
	assign fresh_wire_378[ 3 ] = fresh_wire_878[ 3 ];
	assign fresh_wire_378[ 4 ] = fresh_wire_878[ 4 ];
	assign fresh_wire_378[ 5 ] = fresh_wire_878[ 5 ];
	assign fresh_wire_378[ 6 ] = fresh_wire_878[ 6 ];
	assign fresh_wire_378[ 7 ] = fresh_wire_878[ 7 ];
	assign fresh_wire_378[ 8 ] = fresh_wire_878[ 8 ];
	assign fresh_wire_378[ 9 ] = fresh_wire_878[ 9 ];
	assign fresh_wire_378[ 10 ] = fresh_wire_878[ 10 ];
	assign fresh_wire_378[ 11 ] = fresh_wire_878[ 11 ];
	assign fresh_wire_378[ 12 ] = fresh_wire_878[ 12 ];
	assign fresh_wire_378[ 13 ] = fresh_wire_878[ 13 ];
	assign fresh_wire_378[ 14 ] = fresh_wire_878[ 14 ];
	assign fresh_wire_378[ 15 ] = fresh_wire_878[ 15 ];
	assign fresh_wire_380[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_381[ 0 ] = fresh_wire_455[ 0 ];
	assign fresh_wire_383[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_384[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_385[ 0 ] = fresh_wire_451[ 0 ];
	assign fresh_wire_387[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_388[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_389[ 0 ] = fresh_wire_443[ 0 ];
	assign fresh_wire_391[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_392[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_393[ 0 ] = fresh_wire_535[ 0 ];
	assign fresh_wire_395[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_396[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_397[ 0 ] = fresh_wire_511[ 0 ];
	assign fresh_wire_399[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_400[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_401[ 0 ] = fresh_wire_495[ 0 ];
	assign fresh_wire_401[ 1 ] = fresh_wire_495[ 1 ];
	assign fresh_wire_403[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_404[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_405[ 0 ] = fresh_wire_471[ 0 ];
	assign fresh_wire_405[ 1 ] = fresh_wire_471[ 1 ];
	assign fresh_wire_405[ 2 ] = fresh_wire_471[ 2 ];
	assign fresh_wire_405[ 3 ] = fresh_wire_471[ 3 ];
	assign fresh_wire_405[ 4 ] = fresh_wire_471[ 4 ];
	assign fresh_wire_405[ 5 ] = fresh_wire_471[ 5 ];
	assign fresh_wire_405[ 6 ] = fresh_wire_471[ 6 ];
	assign fresh_wire_405[ 7 ] = fresh_wire_471[ 7 ];
	assign fresh_wire_405[ 8 ] = fresh_wire_471[ 8 ];
	assign fresh_wire_405[ 9 ] = fresh_wire_471[ 9 ];
	assign fresh_wire_405[ 10 ] = fresh_wire_471[ 10 ];
	assign fresh_wire_405[ 11 ] = fresh_wire_471[ 11 ];
	assign fresh_wire_405[ 12 ] = fresh_wire_471[ 12 ];
	assign fresh_wire_405[ 13 ] = fresh_wire_471[ 13 ];
	assign fresh_wire_405[ 14 ] = fresh_wire_471[ 14 ];
	assign fresh_wire_405[ 15 ] = fresh_wire_471[ 15 ];
	assign fresh_wire_407[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_408[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_409[ 0 ] = fresh_wire_571[ 0 ];
	assign fresh_wire_409[ 1 ] = fresh_wire_571[ 1 ];
	assign fresh_wire_409[ 2 ] = fresh_wire_571[ 2 ];
	assign fresh_wire_409[ 3 ] = fresh_wire_571[ 3 ];
	assign fresh_wire_409[ 4 ] = fresh_wire_571[ 4 ];
	assign fresh_wire_409[ 5 ] = fresh_wire_571[ 5 ];
	assign fresh_wire_409[ 6 ] = fresh_wire_571[ 6 ];
	assign fresh_wire_409[ 7 ] = fresh_wire_571[ 7 ];
	assign fresh_wire_409[ 8 ] = fresh_wire_571[ 8 ];
	assign fresh_wire_409[ 9 ] = fresh_wire_571[ 9 ];
	assign fresh_wire_409[ 10 ] = fresh_wire_571[ 10 ];
	assign fresh_wire_409[ 11 ] = fresh_wire_571[ 11 ];
	assign fresh_wire_409[ 12 ] = fresh_wire_571[ 12 ];
	assign fresh_wire_409[ 13 ] = fresh_wire_571[ 13 ];
	assign fresh_wire_409[ 14 ] = fresh_wire_571[ 14 ];
	assign fresh_wire_409[ 15 ] = fresh_wire_571[ 15 ];
	assign fresh_wire_411[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_412[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_413[ 0 ] = fresh_wire_559[ 0 ];
	assign fresh_wire_413[ 1 ] = fresh_wire_559[ 1 ];
	assign fresh_wire_413[ 2 ] = fresh_wire_559[ 2 ];
	assign fresh_wire_413[ 3 ] = fresh_wire_559[ 3 ];
	assign fresh_wire_413[ 4 ] = fresh_wire_559[ 4 ];
	assign fresh_wire_413[ 5 ] = fresh_wire_559[ 5 ];
	assign fresh_wire_413[ 6 ] = fresh_wire_559[ 6 ];
	assign fresh_wire_413[ 7 ] = fresh_wire_559[ 7 ];
	assign fresh_wire_413[ 8 ] = fresh_wire_559[ 8 ];
	assign fresh_wire_413[ 9 ] = fresh_wire_559[ 9 ];
	assign fresh_wire_413[ 10 ] = fresh_wire_559[ 10 ];
	assign fresh_wire_413[ 11 ] = fresh_wire_559[ 11 ];
	assign fresh_wire_413[ 12 ] = fresh_wire_559[ 12 ];
	assign fresh_wire_413[ 13 ] = fresh_wire_559[ 13 ];
	assign fresh_wire_413[ 14 ] = fresh_wire_559[ 14 ];
	assign fresh_wire_413[ 15 ] = fresh_wire_559[ 15 ];
	assign fresh_wire_415[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_416[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_417[ 0 ] = fresh_wire_547[ 0 ];
	assign fresh_wire_417[ 1 ] = fresh_wire_547[ 1 ];
	assign fresh_wire_417[ 2 ] = fresh_wire_547[ 2 ];
	assign fresh_wire_417[ 3 ] = fresh_wire_547[ 3 ];
	assign fresh_wire_417[ 4 ] = fresh_wire_547[ 4 ];
	assign fresh_wire_417[ 5 ] = fresh_wire_547[ 5 ];
	assign fresh_wire_417[ 6 ] = fresh_wire_547[ 6 ];
	assign fresh_wire_417[ 7 ] = fresh_wire_547[ 7 ];
	assign fresh_wire_417[ 8 ] = fresh_wire_547[ 8 ];
	assign fresh_wire_417[ 9 ] = fresh_wire_547[ 9 ];
	assign fresh_wire_417[ 10 ] = fresh_wire_547[ 10 ];
	assign fresh_wire_417[ 11 ] = fresh_wire_547[ 11 ];
	assign fresh_wire_417[ 12 ] = fresh_wire_547[ 12 ];
	assign fresh_wire_417[ 13 ] = fresh_wire_547[ 13 ];
	assign fresh_wire_417[ 14 ] = fresh_wire_547[ 14 ];
	assign fresh_wire_417[ 15 ] = fresh_wire_547[ 15 ];
	assign fresh_wire_419[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_420[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_421[ 0 ] = fresh_wire_591[ 0 ];
	assign fresh_wire_423[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_424[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_425[ 0 ] = fresh_wire_579[ 0 ];
	assign fresh_wire_427[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_428[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_429[ 0 ] = fresh_wire_368[ 0 ];
	assign fresh_wire_431[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_432[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_433[ 0 ] = fresh_wire_414[ 0 ];
	assign fresh_wire_433[ 1 ] = fresh_wire_414[ 1 ];
	assign fresh_wire_433[ 2 ] = fresh_wire_414[ 2 ];
	assign fresh_wire_433[ 3 ] = fresh_wire_414[ 3 ];
	assign fresh_wire_433[ 4 ] = fresh_wire_414[ 4 ];
	assign fresh_wire_433[ 5 ] = fresh_wire_414[ 5 ];
	assign fresh_wire_433[ 6 ] = fresh_wire_414[ 6 ];
	assign fresh_wire_433[ 7 ] = fresh_wire_414[ 7 ];
	assign fresh_wire_433[ 8 ] = fresh_wire_414[ 8 ];
	assign fresh_wire_433[ 9 ] = fresh_wire_414[ 9 ];
	assign fresh_wire_433[ 10 ] = fresh_wire_414[ 10 ];
	assign fresh_wire_433[ 11 ] = fresh_wire_414[ 11 ];
	assign fresh_wire_433[ 12 ] = fresh_wire_414[ 12 ];
	assign fresh_wire_433[ 13 ] = fresh_wire_414[ 13 ];
	assign fresh_wire_433[ 14 ] = fresh_wire_414[ 14 ];
	assign fresh_wire_433[ 15 ] = fresh_wire_414[ 15 ];
	assign fresh_wire_434[ 0 ] = fresh_wire_410[ 0 ];
	assign fresh_wire_434[ 1 ] = fresh_wire_410[ 1 ];
	assign fresh_wire_434[ 2 ] = fresh_wire_410[ 2 ];
	assign fresh_wire_434[ 3 ] = fresh_wire_410[ 3 ];
	assign fresh_wire_434[ 4 ] = fresh_wire_410[ 4 ];
	assign fresh_wire_434[ 5 ] = fresh_wire_410[ 5 ];
	assign fresh_wire_434[ 6 ] = fresh_wire_410[ 6 ];
	assign fresh_wire_434[ 7 ] = fresh_wire_410[ 7 ];
	assign fresh_wire_434[ 8 ] = fresh_wire_410[ 8 ];
	assign fresh_wire_434[ 9 ] = fresh_wire_410[ 9 ];
	assign fresh_wire_434[ 10 ] = fresh_wire_410[ 10 ];
	assign fresh_wire_434[ 11 ] = fresh_wire_410[ 11 ];
	assign fresh_wire_434[ 12 ] = fresh_wire_410[ 12 ];
	assign fresh_wire_434[ 13 ] = fresh_wire_410[ 13 ];
	assign fresh_wire_434[ 14 ] = fresh_wire_410[ 14 ];
	assign fresh_wire_434[ 15 ] = fresh_wire_410[ 15 ];
	assign fresh_wire_436[ 0 ] = fresh_wire_219[ 0 ];
	assign fresh_wire_437[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_438[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_440[ 0 ] = fresh_wire_249[ 0 ];
	assign fresh_wire_441[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_442[ 0 ] = fresh_wire_439[ 0 ];
	assign fresh_wire_444[ 0 ] = fresh_wire_219[ 0 ];
	assign fresh_wire_445[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_446[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_448[ 0 ] = fresh_wire_348[ 0 ];
	assign fresh_wire_449[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_450[ 0 ] = fresh_wire_447[ 0 ];
	assign fresh_wire_452[ 0 ] = fresh_wire_219[ 0 ];
	assign fresh_wire_453[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_454[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_456[ 0 ] = fresh_wire_355[ 0 ];
	assign fresh_wire_457[ 0 ] = fresh_wire_406[ 0 ];
	assign fresh_wire_457[ 1 ] = fresh_wire_406[ 1 ];
	assign fresh_wire_457[ 2 ] = fresh_wire_406[ 2 ];
	assign fresh_wire_457[ 3 ] = fresh_wire_406[ 3 ];
	assign fresh_wire_457[ 4 ] = fresh_wire_406[ 4 ];
	assign fresh_wire_457[ 5 ] = fresh_wire_406[ 5 ];
	assign fresh_wire_457[ 6 ] = fresh_wire_406[ 6 ];
	assign fresh_wire_457[ 7 ] = fresh_wire_406[ 7 ];
	assign fresh_wire_457[ 8 ] = fresh_wire_406[ 8 ];
	assign fresh_wire_457[ 9 ] = fresh_wire_406[ 9 ];
	assign fresh_wire_457[ 10 ] = fresh_wire_406[ 10 ];
	assign fresh_wire_457[ 11 ] = fresh_wire_406[ 11 ];
	assign fresh_wire_457[ 12 ] = fresh_wire_406[ 12 ];
	assign fresh_wire_457[ 13 ] = fresh_wire_406[ 13 ];
	assign fresh_wire_457[ 14 ] = fresh_wire_406[ 14 ];
	assign fresh_wire_457[ 15 ] = fresh_wire_406[ 15 ];
	assign fresh_wire_458[ 0 ] = fresh_wire_192[ 0 ];
	assign fresh_wire_458[ 1 ] = fresh_wire_192[ 1 ];
	assign fresh_wire_458[ 2 ] = fresh_wire_192[ 2 ];
	assign fresh_wire_458[ 3 ] = fresh_wire_192[ 3 ];
	assign fresh_wire_458[ 4 ] = fresh_wire_192[ 4 ];
	assign fresh_wire_458[ 5 ] = fresh_wire_192[ 5 ];
	assign fresh_wire_458[ 6 ] = fresh_wire_192[ 6 ];
	assign fresh_wire_458[ 7 ] = fresh_wire_192[ 7 ];
	assign fresh_wire_458[ 8 ] = fresh_wire_192[ 8 ];
	assign fresh_wire_458[ 9 ] = fresh_wire_192[ 9 ];
	assign fresh_wire_458[ 10 ] = fresh_wire_192[ 10 ];
	assign fresh_wire_458[ 11 ] = fresh_wire_192[ 11 ];
	assign fresh_wire_458[ 12 ] = fresh_wire_192[ 12 ];
	assign fresh_wire_458[ 13 ] = fresh_wire_192[ 13 ];
	assign fresh_wire_458[ 14 ] = fresh_wire_192[ 14 ];
	assign fresh_wire_458[ 15 ] = fresh_wire_192[ 15 ];
	assign fresh_wire_460[ 0 ] = fresh_wire_317[ 0 ];
	assign fresh_wire_461[ 0 ] = fresh_wire_459[ 0 ];
	assign fresh_wire_461[ 1 ] = fresh_wire_459[ 1 ];
	assign fresh_wire_461[ 2 ] = fresh_wire_459[ 2 ];
	assign fresh_wire_461[ 3 ] = fresh_wire_459[ 3 ];
	assign fresh_wire_461[ 4 ] = fresh_wire_459[ 4 ];
	assign fresh_wire_461[ 5 ] = fresh_wire_459[ 5 ];
	assign fresh_wire_461[ 6 ] = fresh_wire_459[ 6 ];
	assign fresh_wire_461[ 7 ] = fresh_wire_459[ 7 ];
	assign fresh_wire_461[ 8 ] = fresh_wire_459[ 8 ];
	assign fresh_wire_461[ 9 ] = fresh_wire_459[ 9 ];
	assign fresh_wire_461[ 10 ] = fresh_wire_459[ 10 ];
	assign fresh_wire_461[ 11 ] = fresh_wire_459[ 11 ];
	assign fresh_wire_461[ 12 ] = fresh_wire_459[ 12 ];
	assign fresh_wire_461[ 13 ] = fresh_wire_459[ 13 ];
	assign fresh_wire_461[ 14 ] = fresh_wire_459[ 14 ];
	assign fresh_wire_461[ 15 ] = fresh_wire_459[ 15 ];
	assign fresh_wire_462[ 0 ] = fresh_wire_604[ 0 ];
	assign fresh_wire_462[ 1 ] = fresh_wire_604[ 1 ];
	assign fresh_wire_462[ 2 ] = fresh_wire_604[ 2 ];
	assign fresh_wire_462[ 3 ] = fresh_wire_604[ 3 ];
	assign fresh_wire_462[ 4 ] = fresh_wire_604[ 4 ];
	assign fresh_wire_462[ 5 ] = fresh_wire_604[ 5 ];
	assign fresh_wire_462[ 6 ] = fresh_wire_604[ 6 ];
	assign fresh_wire_462[ 7 ] = fresh_wire_604[ 7 ];
	assign fresh_wire_462[ 8 ] = fresh_wire_604[ 8 ];
	assign fresh_wire_462[ 9 ] = fresh_wire_604[ 9 ];
	assign fresh_wire_462[ 10 ] = fresh_wire_604[ 10 ];
	assign fresh_wire_462[ 11 ] = fresh_wire_604[ 11 ];
	assign fresh_wire_462[ 12 ] = fresh_wire_604[ 12 ];
	assign fresh_wire_462[ 13 ] = fresh_wire_604[ 13 ];
	assign fresh_wire_462[ 14 ] = fresh_wire_604[ 14 ];
	assign fresh_wire_462[ 15 ] = fresh_wire_604[ 15 ];
	assign fresh_wire_464[ 0 ] = fresh_wire_310[ 0 ];
	assign fresh_wire_465[ 0 ] = fresh_wire_463[ 0 ];
	assign fresh_wire_465[ 1 ] = fresh_wire_463[ 1 ];
	assign fresh_wire_465[ 2 ] = fresh_wire_463[ 2 ];
	assign fresh_wire_465[ 3 ] = fresh_wire_463[ 3 ];
	assign fresh_wire_465[ 4 ] = fresh_wire_463[ 4 ];
	assign fresh_wire_465[ 5 ] = fresh_wire_463[ 5 ];
	assign fresh_wire_465[ 6 ] = fresh_wire_463[ 6 ];
	assign fresh_wire_465[ 7 ] = fresh_wire_463[ 7 ];
	assign fresh_wire_465[ 8 ] = fresh_wire_463[ 8 ];
	assign fresh_wire_465[ 9 ] = fresh_wire_463[ 9 ];
	assign fresh_wire_465[ 10 ] = fresh_wire_463[ 10 ];
	assign fresh_wire_465[ 11 ] = fresh_wire_463[ 11 ];
	assign fresh_wire_465[ 12 ] = fresh_wire_463[ 12 ];
	assign fresh_wire_465[ 13 ] = fresh_wire_463[ 13 ];
	assign fresh_wire_465[ 14 ] = fresh_wire_463[ 14 ];
	assign fresh_wire_465[ 15 ] = fresh_wire_463[ 15 ];
	assign fresh_wire_466[ 0 ] = fresh_wire_406[ 0 ];
	assign fresh_wire_466[ 1 ] = fresh_wire_406[ 1 ];
	assign fresh_wire_466[ 2 ] = fresh_wire_406[ 2 ];
	assign fresh_wire_466[ 3 ] = fresh_wire_406[ 3 ];
	assign fresh_wire_466[ 4 ] = fresh_wire_406[ 4 ];
	assign fresh_wire_466[ 5 ] = fresh_wire_406[ 5 ];
	assign fresh_wire_466[ 6 ] = fresh_wire_406[ 6 ];
	assign fresh_wire_466[ 7 ] = fresh_wire_406[ 7 ];
	assign fresh_wire_466[ 8 ] = fresh_wire_406[ 8 ];
	assign fresh_wire_466[ 9 ] = fresh_wire_406[ 9 ];
	assign fresh_wire_466[ 10 ] = fresh_wire_406[ 10 ];
	assign fresh_wire_466[ 11 ] = fresh_wire_406[ 11 ];
	assign fresh_wire_466[ 12 ] = fresh_wire_406[ 12 ];
	assign fresh_wire_466[ 13 ] = fresh_wire_406[ 13 ];
	assign fresh_wire_466[ 14 ] = fresh_wire_406[ 14 ];
	assign fresh_wire_466[ 15 ] = fresh_wire_406[ 15 ];
	assign fresh_wire_468[ 0 ] = fresh_wire_298[ 0 ];
	assign fresh_wire_469[ 0 ] = fresh_wire_406[ 0 ];
	assign fresh_wire_469[ 1 ] = fresh_wire_406[ 1 ];
	assign fresh_wire_469[ 2 ] = fresh_wire_406[ 2 ];
	assign fresh_wire_469[ 3 ] = fresh_wire_406[ 3 ];
	assign fresh_wire_469[ 4 ] = fresh_wire_406[ 4 ];
	assign fresh_wire_469[ 5 ] = fresh_wire_406[ 5 ];
	assign fresh_wire_469[ 6 ] = fresh_wire_406[ 6 ];
	assign fresh_wire_469[ 7 ] = fresh_wire_406[ 7 ];
	assign fresh_wire_469[ 8 ] = fresh_wire_406[ 8 ];
	assign fresh_wire_469[ 9 ] = fresh_wire_406[ 9 ];
	assign fresh_wire_469[ 10 ] = fresh_wire_406[ 10 ];
	assign fresh_wire_469[ 11 ] = fresh_wire_406[ 11 ];
	assign fresh_wire_469[ 12 ] = fresh_wire_406[ 12 ];
	assign fresh_wire_469[ 13 ] = fresh_wire_406[ 13 ];
	assign fresh_wire_469[ 14 ] = fresh_wire_406[ 14 ];
	assign fresh_wire_469[ 15 ] = fresh_wire_406[ 15 ];
	assign fresh_wire_470[ 0 ] = fresh_wire_467[ 0 ];
	assign fresh_wire_470[ 1 ] = fresh_wire_467[ 1 ];
	assign fresh_wire_470[ 2 ] = fresh_wire_467[ 2 ];
	assign fresh_wire_470[ 3 ] = fresh_wire_467[ 3 ];
	assign fresh_wire_470[ 4 ] = fresh_wire_467[ 4 ];
	assign fresh_wire_470[ 5 ] = fresh_wire_467[ 5 ];
	assign fresh_wire_470[ 6 ] = fresh_wire_467[ 6 ];
	assign fresh_wire_470[ 7 ] = fresh_wire_467[ 7 ];
	assign fresh_wire_470[ 8 ] = fresh_wire_467[ 8 ];
	assign fresh_wire_470[ 9 ] = fresh_wire_467[ 9 ];
	assign fresh_wire_470[ 10 ] = fresh_wire_467[ 10 ];
	assign fresh_wire_470[ 11 ] = fresh_wire_467[ 11 ];
	assign fresh_wire_470[ 12 ] = fresh_wire_467[ 12 ];
	assign fresh_wire_470[ 13 ] = fresh_wire_467[ 13 ];
	assign fresh_wire_470[ 14 ] = fresh_wire_467[ 14 ];
	assign fresh_wire_470[ 15 ] = fresh_wire_467[ 15 ];
	assign fresh_wire_472[ 0 ] = fresh_wire_219[ 0 ];
	assign fresh_wire_473[ 0 ] = fresh_wire_402[ 0 ];
	assign fresh_wire_473[ 1 ] = fresh_wire_402[ 1 ];
	assign fresh_wire_474[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_474[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_476[ 0 ] = fresh_wire_329[ 0 ];
	assign fresh_wire_477[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_477[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_478[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_478[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_480[ 0 ] = fresh_wire_322[ 0 ];
	assign fresh_wire_481[ 0 ] = fresh_wire_475[ 0 ];
	assign fresh_wire_481[ 1 ] = fresh_wire_475[ 1 ];
	assign fresh_wire_482[ 0 ] = fresh_wire_479[ 0 ];
	assign fresh_wire_482[ 1 ] = fresh_wire_479[ 1 ];
	assign fresh_wire_484[ 0 ] = fresh_wire_317[ 0 ];
	assign fresh_wire_485[ 0 ] = fresh_wire_483[ 0 ];
	assign fresh_wire_485[ 1 ] = fresh_wire_483[ 1 ];
	assign fresh_wire_486[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_486[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_488[ 0 ] = fresh_wire_310[ 0 ];
	assign fresh_wire_489[ 0 ] = fresh_wire_487[ 0 ];
	assign fresh_wire_489[ 1 ] = fresh_wire_487[ 1 ];
	assign fresh_wire_490[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_490[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_492[ 0 ] = fresh_wire_298[ 0 ];
	assign fresh_wire_493[ 0 ] = fresh_wire_402[ 0 ];
	assign fresh_wire_493[ 1 ] = fresh_wire_402[ 1 ];
	assign fresh_wire_494[ 0 ] = fresh_wire_491[ 0 ];
	assign fresh_wire_494[ 1 ] = fresh_wire_491[ 1 ];
	assign fresh_wire_496[ 0 ] = fresh_wire_219[ 0 ];
	assign fresh_wire_497[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_498[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_500[ 0 ] = fresh_wire_317[ 0 ];
	assign fresh_wire_501[ 0 ] = fresh_wire_499[ 0 ];
	assign fresh_wire_502[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_504[ 0 ] = fresh_wire_310[ 0 ];
	assign fresh_wire_505[ 0 ] = fresh_wire_503[ 0 ];
	assign fresh_wire_506[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_508[ 0 ] = fresh_wire_298[ 0 ];
	assign fresh_wire_509[ 0 ] = fresh_wire_398[ 0 ];
	assign fresh_wire_510[ 0 ] = fresh_wire_507[ 0 ];
	assign fresh_wire_512[ 0 ] = fresh_wire_219[ 0 ];
	assign fresh_wire_513[ 0 ] = fresh_wire_394[ 0 ];
	assign fresh_wire_514[ 0 ] = fresh_wire_370[ 0 ];
	assign fresh_wire_516[ 0 ] = fresh_wire_329[ 0 ];
	assign fresh_wire_517[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_518[ 0 ] = fresh_wire_394[ 0 ];
	assign fresh_wire_520[ 0 ] = fresh_wire_322[ 0 ];
	assign fresh_wire_521[ 0 ] = fresh_wire_515[ 0 ];
	assign fresh_wire_522[ 0 ] = fresh_wire_519[ 0 ];
	assign fresh_wire_524[ 0 ] = fresh_wire_317[ 0 ];
	assign fresh_wire_525[ 0 ] = fresh_wire_523[ 0 ];
	assign fresh_wire_526[ 0 ] = fresh_wire_394[ 0 ];
	assign fresh_wire_528[ 0 ] = fresh_wire_310[ 0 ];
	assign fresh_wire_529[ 0 ] = fresh_wire_527[ 0 ];
	assign fresh_wire_530[ 0 ] = fresh_wire_370[ 0 ];
	assign fresh_wire_532[ 0 ] = fresh_wire_298[ 0 ];
	assign fresh_wire_533[ 0 ] = fresh_wire_394[ 0 ];
	assign fresh_wire_534[ 0 ] = fresh_wire_531[ 0 ];
	assign fresh_wire_536[ 0 ] = fresh_wire_219[ 0 ];
	assign fresh_wire_537[ 0 ] = fresh_wire_418[ 0 ];
	assign fresh_wire_537[ 1 ] = fresh_wire_418[ 1 ];
	assign fresh_wire_537[ 2 ] = fresh_wire_418[ 2 ];
	assign fresh_wire_537[ 3 ] = fresh_wire_418[ 3 ];
	assign fresh_wire_537[ 4 ] = fresh_wire_418[ 4 ];
	assign fresh_wire_537[ 5 ] = fresh_wire_418[ 5 ];
	assign fresh_wire_537[ 6 ] = fresh_wire_418[ 6 ];
	assign fresh_wire_537[ 7 ] = fresh_wire_418[ 7 ];
	assign fresh_wire_537[ 8 ] = fresh_wire_418[ 8 ];
	assign fresh_wire_537[ 9 ] = fresh_wire_418[ 9 ];
	assign fresh_wire_537[ 10 ] = fresh_wire_418[ 10 ];
	assign fresh_wire_537[ 11 ] = fresh_wire_418[ 11 ];
	assign fresh_wire_537[ 12 ] = fresh_wire_418[ 12 ];
	assign fresh_wire_537[ 13 ] = fresh_wire_418[ 13 ];
	assign fresh_wire_537[ 14 ] = fresh_wire_418[ 14 ];
	assign fresh_wire_537[ 15 ] = fresh_wire_418[ 15 ];
	assign fresh_wire_538[ 0 ] = fresh_wire_597[ 0 ];
	assign fresh_wire_538[ 1 ] = fresh_wire_597[ 1 ];
	assign fresh_wire_538[ 2 ] = fresh_wire_597[ 2 ];
	assign fresh_wire_538[ 3 ] = fresh_wire_597[ 3 ];
	assign fresh_wire_538[ 4 ] = fresh_wire_597[ 4 ];
	assign fresh_wire_538[ 5 ] = fresh_wire_597[ 5 ];
	assign fresh_wire_538[ 6 ] = fresh_wire_597[ 6 ];
	assign fresh_wire_538[ 7 ] = fresh_wire_597[ 7 ];
	assign fresh_wire_538[ 8 ] = fresh_wire_597[ 8 ];
	assign fresh_wire_538[ 9 ] = fresh_wire_597[ 9 ];
	assign fresh_wire_538[ 10 ] = fresh_wire_597[ 10 ];
	assign fresh_wire_538[ 11 ] = fresh_wire_597[ 11 ];
	assign fresh_wire_538[ 12 ] = fresh_wire_597[ 12 ];
	assign fresh_wire_538[ 13 ] = fresh_wire_597[ 13 ];
	assign fresh_wire_538[ 14 ] = fresh_wire_597[ 14 ];
	assign fresh_wire_538[ 15 ] = fresh_wire_597[ 15 ];
	assign fresh_wire_540[ 0 ] = fresh_wire_228[ 0 ];
	assign fresh_wire_541[ 0 ] = fresh_wire_418[ 0 ];
	assign fresh_wire_541[ 1 ] = fresh_wire_418[ 1 ];
	assign fresh_wire_541[ 2 ] = fresh_wire_418[ 2 ];
	assign fresh_wire_541[ 3 ] = fresh_wire_418[ 3 ];
	assign fresh_wire_541[ 4 ] = fresh_wire_418[ 4 ];
	assign fresh_wire_541[ 5 ] = fresh_wire_418[ 5 ];
	assign fresh_wire_541[ 6 ] = fresh_wire_418[ 6 ];
	assign fresh_wire_541[ 7 ] = fresh_wire_418[ 7 ];
	assign fresh_wire_541[ 8 ] = fresh_wire_418[ 8 ];
	assign fresh_wire_541[ 9 ] = fresh_wire_418[ 9 ];
	assign fresh_wire_541[ 10 ] = fresh_wire_418[ 10 ];
	assign fresh_wire_541[ 11 ] = fresh_wire_418[ 11 ];
	assign fresh_wire_541[ 12 ] = fresh_wire_418[ 12 ];
	assign fresh_wire_541[ 13 ] = fresh_wire_418[ 13 ];
	assign fresh_wire_541[ 14 ] = fresh_wire_418[ 14 ];
	assign fresh_wire_541[ 15 ] = fresh_wire_418[ 15 ];
	assign fresh_wire_542[ 0 ] = fresh_wire_181[ 0 ];
	assign fresh_wire_542[ 1 ] = fresh_wire_181[ 1 ];
	assign fresh_wire_542[ 2 ] = fresh_wire_181[ 2 ];
	assign fresh_wire_542[ 3 ] = fresh_wire_181[ 3 ];
	assign fresh_wire_542[ 4 ] = fresh_wire_181[ 4 ];
	assign fresh_wire_542[ 5 ] = fresh_wire_181[ 5 ];
	assign fresh_wire_542[ 6 ] = fresh_wire_181[ 6 ];
	assign fresh_wire_542[ 7 ] = fresh_wire_181[ 7 ];
	assign fresh_wire_542[ 8 ] = fresh_wire_181[ 8 ];
	assign fresh_wire_542[ 9 ] = fresh_wire_181[ 9 ];
	assign fresh_wire_542[ 10 ] = fresh_wire_181[ 10 ];
	assign fresh_wire_542[ 11 ] = fresh_wire_181[ 11 ];
	assign fresh_wire_542[ 12 ] = fresh_wire_181[ 12 ];
	assign fresh_wire_542[ 13 ] = fresh_wire_181[ 13 ];
	assign fresh_wire_542[ 14 ] = fresh_wire_181[ 14 ];
	assign fresh_wire_542[ 15 ] = fresh_wire_181[ 15 ];
	assign fresh_wire_544[ 0 ] = fresh_wire_234[ 0 ];
	assign fresh_wire_545[ 0 ] = fresh_wire_539[ 0 ];
	assign fresh_wire_545[ 1 ] = fresh_wire_539[ 1 ];
	assign fresh_wire_545[ 2 ] = fresh_wire_539[ 2 ];
	assign fresh_wire_545[ 3 ] = fresh_wire_539[ 3 ];
	assign fresh_wire_545[ 4 ] = fresh_wire_539[ 4 ];
	assign fresh_wire_545[ 5 ] = fresh_wire_539[ 5 ];
	assign fresh_wire_545[ 6 ] = fresh_wire_539[ 6 ];
	assign fresh_wire_545[ 7 ] = fresh_wire_539[ 7 ];
	assign fresh_wire_545[ 8 ] = fresh_wire_539[ 8 ];
	assign fresh_wire_545[ 9 ] = fresh_wire_539[ 9 ];
	assign fresh_wire_545[ 10 ] = fresh_wire_539[ 10 ];
	assign fresh_wire_545[ 11 ] = fresh_wire_539[ 11 ];
	assign fresh_wire_545[ 12 ] = fresh_wire_539[ 12 ];
	assign fresh_wire_545[ 13 ] = fresh_wire_539[ 13 ];
	assign fresh_wire_545[ 14 ] = fresh_wire_539[ 14 ];
	assign fresh_wire_545[ 15 ] = fresh_wire_539[ 15 ];
	assign fresh_wire_546[ 0 ] = fresh_wire_543[ 0 ];
	assign fresh_wire_546[ 1 ] = fresh_wire_543[ 1 ];
	assign fresh_wire_546[ 2 ] = fresh_wire_543[ 2 ];
	assign fresh_wire_546[ 3 ] = fresh_wire_543[ 3 ];
	assign fresh_wire_546[ 4 ] = fresh_wire_543[ 4 ];
	assign fresh_wire_546[ 5 ] = fresh_wire_543[ 5 ];
	assign fresh_wire_546[ 6 ] = fresh_wire_543[ 6 ];
	assign fresh_wire_546[ 7 ] = fresh_wire_543[ 7 ];
	assign fresh_wire_546[ 8 ] = fresh_wire_543[ 8 ];
	assign fresh_wire_546[ 9 ] = fresh_wire_543[ 9 ];
	assign fresh_wire_546[ 10 ] = fresh_wire_543[ 10 ];
	assign fresh_wire_546[ 11 ] = fresh_wire_543[ 11 ];
	assign fresh_wire_546[ 12 ] = fresh_wire_543[ 12 ];
	assign fresh_wire_546[ 13 ] = fresh_wire_543[ 13 ];
	assign fresh_wire_546[ 14 ] = fresh_wire_543[ 14 ];
	assign fresh_wire_546[ 15 ] = fresh_wire_543[ 15 ];
	assign fresh_wire_548[ 0 ] = fresh_wire_231[ 0 ];
	assign fresh_wire_549[ 0 ] = fresh_wire_176[ 0 ];
	assign fresh_wire_549[ 1 ] = fresh_wire_176[ 1 ];
	assign fresh_wire_549[ 2 ] = fresh_wire_176[ 2 ];
	assign fresh_wire_549[ 3 ] = fresh_wire_176[ 3 ];
	assign fresh_wire_549[ 4 ] = fresh_wire_176[ 4 ];
	assign fresh_wire_549[ 5 ] = fresh_wire_176[ 5 ];
	assign fresh_wire_549[ 6 ] = fresh_wire_176[ 6 ];
	assign fresh_wire_549[ 7 ] = fresh_wire_176[ 7 ];
	assign fresh_wire_549[ 8 ] = fresh_wire_176[ 8 ];
	assign fresh_wire_549[ 9 ] = fresh_wire_176[ 9 ];
	assign fresh_wire_549[ 10 ] = fresh_wire_176[ 10 ];
	assign fresh_wire_549[ 11 ] = fresh_wire_176[ 11 ];
	assign fresh_wire_549[ 12 ] = fresh_wire_176[ 12 ];
	assign fresh_wire_549[ 13 ] = fresh_wire_176[ 13 ];
	assign fresh_wire_549[ 14 ] = fresh_wire_176[ 14 ];
	assign fresh_wire_549[ 15 ] = fresh_wire_176[ 15 ];
	assign fresh_wire_550[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_550[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_550[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_550[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_550[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_550[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_550[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_550[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_550[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_550[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_550[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_550[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_550[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_550[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_550[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_550[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_552[ 0 ] = fresh_wire_261[ 0 ];
	assign fresh_wire_553[ 0 ] = fresh_wire_414[ 0 ];
	assign fresh_wire_553[ 1 ] = fresh_wire_414[ 1 ];
	assign fresh_wire_553[ 2 ] = fresh_wire_414[ 2 ];
	assign fresh_wire_553[ 3 ] = fresh_wire_414[ 3 ];
	assign fresh_wire_553[ 4 ] = fresh_wire_414[ 4 ];
	assign fresh_wire_553[ 5 ] = fresh_wire_414[ 5 ];
	assign fresh_wire_553[ 6 ] = fresh_wire_414[ 6 ];
	assign fresh_wire_553[ 7 ] = fresh_wire_414[ 7 ];
	assign fresh_wire_553[ 8 ] = fresh_wire_414[ 8 ];
	assign fresh_wire_553[ 9 ] = fresh_wire_414[ 9 ];
	assign fresh_wire_553[ 10 ] = fresh_wire_414[ 10 ];
	assign fresh_wire_553[ 11 ] = fresh_wire_414[ 11 ];
	assign fresh_wire_553[ 12 ] = fresh_wire_414[ 12 ];
	assign fresh_wire_553[ 13 ] = fresh_wire_414[ 13 ];
	assign fresh_wire_553[ 14 ] = fresh_wire_414[ 14 ];
	assign fresh_wire_553[ 15 ] = fresh_wire_414[ 15 ];
	assign fresh_wire_554[ 0 ] = fresh_wire_551[ 0 ];
	assign fresh_wire_554[ 1 ] = fresh_wire_551[ 1 ];
	assign fresh_wire_554[ 2 ] = fresh_wire_551[ 2 ];
	assign fresh_wire_554[ 3 ] = fresh_wire_551[ 3 ];
	assign fresh_wire_554[ 4 ] = fresh_wire_551[ 4 ];
	assign fresh_wire_554[ 5 ] = fresh_wire_551[ 5 ];
	assign fresh_wire_554[ 6 ] = fresh_wire_551[ 6 ];
	assign fresh_wire_554[ 7 ] = fresh_wire_551[ 7 ];
	assign fresh_wire_554[ 8 ] = fresh_wire_551[ 8 ];
	assign fresh_wire_554[ 9 ] = fresh_wire_551[ 9 ];
	assign fresh_wire_554[ 10 ] = fresh_wire_551[ 10 ];
	assign fresh_wire_554[ 11 ] = fresh_wire_551[ 11 ];
	assign fresh_wire_554[ 12 ] = fresh_wire_551[ 12 ];
	assign fresh_wire_554[ 13 ] = fresh_wire_551[ 13 ];
	assign fresh_wire_554[ 14 ] = fresh_wire_551[ 14 ];
	assign fresh_wire_554[ 15 ] = fresh_wire_551[ 15 ];
	assign fresh_wire_556[ 0 ] = fresh_wire_234[ 0 ];
	assign fresh_wire_557[ 0 ] = fresh_wire_414[ 0 ];
	assign fresh_wire_557[ 1 ] = fresh_wire_414[ 1 ];
	assign fresh_wire_557[ 2 ] = fresh_wire_414[ 2 ];
	assign fresh_wire_557[ 3 ] = fresh_wire_414[ 3 ];
	assign fresh_wire_557[ 4 ] = fresh_wire_414[ 4 ];
	assign fresh_wire_557[ 5 ] = fresh_wire_414[ 5 ];
	assign fresh_wire_557[ 6 ] = fresh_wire_414[ 6 ];
	assign fresh_wire_557[ 7 ] = fresh_wire_414[ 7 ];
	assign fresh_wire_557[ 8 ] = fresh_wire_414[ 8 ];
	assign fresh_wire_557[ 9 ] = fresh_wire_414[ 9 ];
	assign fresh_wire_557[ 10 ] = fresh_wire_414[ 10 ];
	assign fresh_wire_557[ 11 ] = fresh_wire_414[ 11 ];
	assign fresh_wire_557[ 12 ] = fresh_wire_414[ 12 ];
	assign fresh_wire_557[ 13 ] = fresh_wire_414[ 13 ];
	assign fresh_wire_557[ 14 ] = fresh_wire_414[ 14 ];
	assign fresh_wire_557[ 15 ] = fresh_wire_414[ 15 ];
	assign fresh_wire_558[ 0 ] = fresh_wire_555[ 0 ];
	assign fresh_wire_558[ 1 ] = fresh_wire_555[ 1 ];
	assign fresh_wire_558[ 2 ] = fresh_wire_555[ 2 ];
	assign fresh_wire_558[ 3 ] = fresh_wire_555[ 3 ];
	assign fresh_wire_558[ 4 ] = fresh_wire_555[ 4 ];
	assign fresh_wire_558[ 5 ] = fresh_wire_555[ 5 ];
	assign fresh_wire_558[ 6 ] = fresh_wire_555[ 6 ];
	assign fresh_wire_558[ 7 ] = fresh_wire_555[ 7 ];
	assign fresh_wire_558[ 8 ] = fresh_wire_555[ 8 ];
	assign fresh_wire_558[ 9 ] = fresh_wire_555[ 9 ];
	assign fresh_wire_558[ 10 ] = fresh_wire_555[ 10 ];
	assign fresh_wire_558[ 11 ] = fresh_wire_555[ 11 ];
	assign fresh_wire_558[ 12 ] = fresh_wire_555[ 12 ];
	assign fresh_wire_558[ 13 ] = fresh_wire_555[ 13 ];
	assign fresh_wire_558[ 14 ] = fresh_wire_555[ 14 ];
	assign fresh_wire_558[ 15 ] = fresh_wire_555[ 15 ];
	assign fresh_wire_560[ 0 ] = fresh_wire_231[ 0 ];
	assign fresh_wire_561[ 0 ] = fresh_wire_186[ 0 ];
	assign fresh_wire_561[ 1 ] = fresh_wire_186[ 1 ];
	assign fresh_wire_561[ 2 ] = fresh_wire_186[ 2 ];
	assign fresh_wire_561[ 3 ] = fresh_wire_186[ 3 ];
	assign fresh_wire_561[ 4 ] = fresh_wire_186[ 4 ];
	assign fresh_wire_561[ 5 ] = fresh_wire_186[ 5 ];
	assign fresh_wire_561[ 6 ] = fresh_wire_186[ 6 ];
	assign fresh_wire_561[ 7 ] = fresh_wire_186[ 7 ];
	assign fresh_wire_561[ 8 ] = fresh_wire_186[ 8 ];
	assign fresh_wire_561[ 9 ] = fresh_wire_186[ 9 ];
	assign fresh_wire_561[ 10 ] = fresh_wire_186[ 10 ];
	assign fresh_wire_561[ 11 ] = fresh_wire_186[ 11 ];
	assign fresh_wire_561[ 12 ] = fresh_wire_186[ 12 ];
	assign fresh_wire_561[ 13 ] = fresh_wire_186[ 13 ];
	assign fresh_wire_561[ 14 ] = fresh_wire_186[ 14 ];
	assign fresh_wire_561[ 15 ] = fresh_wire_186[ 15 ];
	assign fresh_wire_562[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_562[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_562[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_562[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_562[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_562[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_562[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_562[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_562[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_562[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_562[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_562[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_562[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_562[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_562[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_562[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_564[ 0 ] = fresh_wire_264[ 0 ];
	assign fresh_wire_565[ 0 ] = fresh_wire_410[ 0 ];
	assign fresh_wire_565[ 1 ] = fresh_wire_410[ 1 ];
	assign fresh_wire_565[ 2 ] = fresh_wire_410[ 2 ];
	assign fresh_wire_565[ 3 ] = fresh_wire_410[ 3 ];
	assign fresh_wire_565[ 4 ] = fresh_wire_410[ 4 ];
	assign fresh_wire_565[ 5 ] = fresh_wire_410[ 5 ];
	assign fresh_wire_565[ 6 ] = fresh_wire_410[ 6 ];
	assign fresh_wire_565[ 7 ] = fresh_wire_410[ 7 ];
	assign fresh_wire_565[ 8 ] = fresh_wire_410[ 8 ];
	assign fresh_wire_565[ 9 ] = fresh_wire_410[ 9 ];
	assign fresh_wire_565[ 10 ] = fresh_wire_410[ 10 ];
	assign fresh_wire_565[ 11 ] = fresh_wire_410[ 11 ];
	assign fresh_wire_565[ 12 ] = fresh_wire_410[ 12 ];
	assign fresh_wire_565[ 13 ] = fresh_wire_410[ 13 ];
	assign fresh_wire_565[ 14 ] = fresh_wire_410[ 14 ];
	assign fresh_wire_565[ 15 ] = fresh_wire_410[ 15 ];
	assign fresh_wire_566[ 0 ] = fresh_wire_563[ 0 ];
	assign fresh_wire_566[ 1 ] = fresh_wire_563[ 1 ];
	assign fresh_wire_566[ 2 ] = fresh_wire_563[ 2 ];
	assign fresh_wire_566[ 3 ] = fresh_wire_563[ 3 ];
	assign fresh_wire_566[ 4 ] = fresh_wire_563[ 4 ];
	assign fresh_wire_566[ 5 ] = fresh_wire_563[ 5 ];
	assign fresh_wire_566[ 6 ] = fresh_wire_563[ 6 ];
	assign fresh_wire_566[ 7 ] = fresh_wire_563[ 7 ];
	assign fresh_wire_566[ 8 ] = fresh_wire_563[ 8 ];
	assign fresh_wire_566[ 9 ] = fresh_wire_563[ 9 ];
	assign fresh_wire_566[ 10 ] = fresh_wire_563[ 10 ];
	assign fresh_wire_566[ 11 ] = fresh_wire_563[ 11 ];
	assign fresh_wire_566[ 12 ] = fresh_wire_563[ 12 ];
	assign fresh_wire_566[ 13 ] = fresh_wire_563[ 13 ];
	assign fresh_wire_566[ 14 ] = fresh_wire_563[ 14 ];
	assign fresh_wire_566[ 15 ] = fresh_wire_563[ 15 ];
	assign fresh_wire_568[ 0 ] = fresh_wire_228[ 0 ];
	assign fresh_wire_569[ 0 ] = fresh_wire_567[ 0 ];
	assign fresh_wire_569[ 1 ] = fresh_wire_567[ 1 ];
	assign fresh_wire_569[ 2 ] = fresh_wire_567[ 2 ];
	assign fresh_wire_569[ 3 ] = fresh_wire_567[ 3 ];
	assign fresh_wire_569[ 4 ] = fresh_wire_567[ 4 ];
	assign fresh_wire_569[ 5 ] = fresh_wire_567[ 5 ];
	assign fresh_wire_569[ 6 ] = fresh_wire_567[ 6 ];
	assign fresh_wire_569[ 7 ] = fresh_wire_567[ 7 ];
	assign fresh_wire_569[ 8 ] = fresh_wire_567[ 8 ];
	assign fresh_wire_569[ 9 ] = fresh_wire_567[ 9 ];
	assign fresh_wire_569[ 10 ] = fresh_wire_567[ 10 ];
	assign fresh_wire_569[ 11 ] = fresh_wire_567[ 11 ];
	assign fresh_wire_569[ 12 ] = fresh_wire_567[ 12 ];
	assign fresh_wire_569[ 13 ] = fresh_wire_567[ 13 ];
	assign fresh_wire_569[ 14 ] = fresh_wire_567[ 14 ];
	assign fresh_wire_569[ 15 ] = fresh_wire_567[ 15 ];
	assign fresh_wire_570[ 0 ] = fresh_wire_410[ 0 ];
	assign fresh_wire_570[ 1 ] = fresh_wire_410[ 1 ];
	assign fresh_wire_570[ 2 ] = fresh_wire_410[ 2 ];
	assign fresh_wire_570[ 3 ] = fresh_wire_410[ 3 ];
	assign fresh_wire_570[ 4 ] = fresh_wire_410[ 4 ];
	assign fresh_wire_570[ 5 ] = fresh_wire_410[ 5 ];
	assign fresh_wire_570[ 6 ] = fresh_wire_410[ 6 ];
	assign fresh_wire_570[ 7 ] = fresh_wire_410[ 7 ];
	assign fresh_wire_570[ 8 ] = fresh_wire_410[ 8 ];
	assign fresh_wire_570[ 9 ] = fresh_wire_410[ 9 ];
	assign fresh_wire_570[ 10 ] = fresh_wire_410[ 10 ];
	assign fresh_wire_570[ 11 ] = fresh_wire_410[ 11 ];
	assign fresh_wire_570[ 12 ] = fresh_wire_410[ 12 ];
	assign fresh_wire_570[ 13 ] = fresh_wire_410[ 13 ];
	assign fresh_wire_570[ 14 ] = fresh_wire_410[ 14 ];
	assign fresh_wire_570[ 15 ] = fresh_wire_410[ 15 ];
	assign fresh_wire_572[ 0 ] = fresh_wire_231[ 0 ];
	assign fresh_wire_573[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_574[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_576[ 0 ] = fresh_wire_222[ 0 ];
	assign fresh_wire_577[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_578[ 0 ] = fresh_wire_575[ 0 ];
	assign fresh_wire_580[ 0 ] = fresh_wire_219[ 0 ];
	assign fresh_wire_581[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_582[ 0 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_584[ 0 ] = fresh_wire_225[ 0 ];
	assign fresh_wire_585[ 0 ] = fresh_wire_583[ 0 ];
	assign fresh_wire_586[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_588[ 0 ] = fresh_wire_222[ 0 ];
	assign fresh_wire_589[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_590[ 0 ] = fresh_wire_587[ 0 ];
	assign fresh_wire_592[ 0 ] = fresh_wire_219[ 0 ];
	assign fresh_wire_593[ 0 ] = fresh_wire_418[ 0 ];
	assign fresh_wire_593[ 1 ] = fresh_wire_418[ 1 ];
	assign fresh_wire_593[ 2 ] = fresh_wire_418[ 2 ];
	assign fresh_wire_593[ 3 ] = fresh_wire_418[ 3 ];
	assign fresh_wire_593[ 4 ] = fresh_wire_418[ 4 ];
	assign fresh_wire_593[ 5 ] = fresh_wire_418[ 5 ];
	assign fresh_wire_593[ 6 ] = fresh_wire_418[ 6 ];
	assign fresh_wire_593[ 7 ] = fresh_wire_418[ 7 ];
	assign fresh_wire_593[ 8 ] = fresh_wire_418[ 8 ];
	assign fresh_wire_593[ 9 ] = fresh_wire_418[ 9 ];
	assign fresh_wire_593[ 10 ] = fresh_wire_418[ 10 ];
	assign fresh_wire_593[ 11 ] = fresh_wire_418[ 11 ];
	assign fresh_wire_593[ 12 ] = fresh_wire_418[ 12 ];
	assign fresh_wire_593[ 13 ] = fresh_wire_418[ 13 ];
	assign fresh_wire_593[ 14 ] = fresh_wire_418[ 14 ];
	assign fresh_wire_593[ 15 ] = fresh_wire_418[ 15 ];
	assign fresh_wire_595[ 0 ] = fresh_wire_594[ 0 ];
	assign fresh_wire_595[ 1 ] = fresh_wire_594[ 1 ];
	assign fresh_wire_595[ 2 ] = fresh_wire_594[ 2 ];
	assign fresh_wire_595[ 3 ] = fresh_wire_594[ 3 ];
	assign fresh_wire_595[ 4 ] = fresh_wire_594[ 4 ];
	assign fresh_wire_595[ 5 ] = fresh_wire_594[ 5 ];
	assign fresh_wire_595[ 6 ] = fresh_wire_594[ 6 ];
	assign fresh_wire_595[ 7 ] = fresh_wire_594[ 7 ];
	assign fresh_wire_595[ 8 ] = fresh_wire_594[ 8 ];
	assign fresh_wire_595[ 9 ] = fresh_wire_594[ 9 ];
	assign fresh_wire_595[ 10 ] = fresh_wire_594[ 10 ];
	assign fresh_wire_595[ 11 ] = fresh_wire_594[ 11 ];
	assign fresh_wire_595[ 12 ] = fresh_wire_594[ 12 ];
	assign fresh_wire_595[ 13 ] = fresh_wire_594[ 13 ];
	assign fresh_wire_595[ 14 ] = fresh_wire_594[ 14 ];
	assign fresh_wire_595[ 15 ] = fresh_wire_594[ 15 ];
	assign fresh_wire_595[ 16 ] = fresh_wire_594[ 16 ];
	assign fresh_wire_595[ 17 ] = fresh_wire_594[ 17 ];
	assign fresh_wire_595[ 18 ] = fresh_wire_594[ 18 ];
	assign fresh_wire_595[ 19 ] = fresh_wire_594[ 19 ];
	assign fresh_wire_595[ 20 ] = fresh_wire_594[ 20 ];
	assign fresh_wire_595[ 21 ] = fresh_wire_594[ 21 ];
	assign fresh_wire_595[ 22 ] = fresh_wire_594[ 22 ];
	assign fresh_wire_595[ 23 ] = fresh_wire_594[ 23 ];
	assign fresh_wire_595[ 24 ] = fresh_wire_594[ 24 ];
	assign fresh_wire_595[ 25 ] = fresh_wire_594[ 25 ];
	assign fresh_wire_595[ 26 ] = fresh_wire_594[ 26 ];
	assign fresh_wire_595[ 27 ] = fresh_wire_594[ 27 ];
	assign fresh_wire_595[ 28 ] = fresh_wire_594[ 28 ];
	assign fresh_wire_595[ 29 ] = fresh_wire_594[ 29 ];
	assign fresh_wire_595[ 30 ] = fresh_wire_594[ 30 ];
	assign fresh_wire_595[ 31 ] = fresh_wire_594[ 31 ];
	assign fresh_wire_596[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 1 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_596[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 16 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 17 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 18 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 19 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 20 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 21 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 22 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 23 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 24 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 25 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 26 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 27 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 28 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 29 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 30 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_596[ 31 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_598[ 0 ] = fresh_wire_939[ 0 ];
	assign fresh_wire_598[ 1 ] = fresh_wire_939[ 1 ];
	assign fresh_wire_598[ 2 ] = fresh_wire_939[ 2 ];
	assign fresh_wire_598[ 3 ] = fresh_wire_939[ 3 ];
	assign fresh_wire_598[ 4 ] = fresh_wire_939[ 4 ];
	assign fresh_wire_598[ 5 ] = fresh_wire_939[ 5 ];
	assign fresh_wire_598[ 6 ] = fresh_wire_939[ 6 ];
	assign fresh_wire_598[ 7 ] = fresh_wire_939[ 7 ];
	assign fresh_wire_598[ 8 ] = fresh_wire_939[ 8 ];
	assign fresh_wire_598[ 9 ] = fresh_wire_939[ 9 ];
	assign fresh_wire_598[ 10 ] = fresh_wire_939[ 10 ];
	assign fresh_wire_598[ 11 ] = fresh_wire_939[ 11 ];
	assign fresh_wire_598[ 12 ] = fresh_wire_939[ 12 ];
	assign fresh_wire_598[ 13 ] = fresh_wire_939[ 13 ];
	assign fresh_wire_598[ 14 ] = fresh_wire_939[ 14 ];
	assign fresh_wire_598[ 15 ] = fresh_wire_939[ 15 ];
	assign fresh_wire_598[ 16 ] = fresh_wire_1037[ 0 ];
	assign fresh_wire_598[ 17 ] = fresh_wire_1037[ 1 ];
	assign fresh_wire_598[ 18 ] = fresh_wire_1037[ 2 ];
	assign fresh_wire_598[ 19 ] = fresh_wire_1037[ 3 ];
	assign fresh_wire_598[ 20 ] = fresh_wire_1037[ 4 ];
	assign fresh_wire_598[ 21 ] = fresh_wire_1037[ 5 ];
	assign fresh_wire_598[ 22 ] = fresh_wire_1037[ 6 ];
	assign fresh_wire_598[ 23 ] = fresh_wire_1037[ 7 ];
	assign fresh_wire_598[ 24 ] = fresh_wire_1037[ 8 ];
	assign fresh_wire_598[ 25 ] = fresh_wire_1037[ 9 ];
	assign fresh_wire_598[ 26 ] = fresh_wire_1037[ 10 ];
	assign fresh_wire_598[ 27 ] = fresh_wire_1037[ 11 ];
	assign fresh_wire_598[ 28 ] = fresh_wire_1037[ 12 ];
	assign fresh_wire_598[ 29 ] = fresh_wire_1037[ 13 ];
	assign fresh_wire_598[ 30 ] = fresh_wire_1037[ 14 ];
	assign fresh_wire_598[ 31 ] = fresh_wire_1037[ 15 ];
	assign fresh_wire_599[ 0 ] = fresh_wire_714[ 0 ];
	assign fresh_wire_599[ 1 ] = fresh_wire_714[ 1 ];
	assign fresh_wire_599[ 2 ] = fresh_wire_714[ 2 ];
	assign fresh_wire_599[ 3 ] = fresh_wire_714[ 3 ];
	assign fresh_wire_599[ 4 ] = fresh_wire_714[ 4 ];
	assign fresh_wire_599[ 5 ] = fresh_wire_714[ 5 ];
	assign fresh_wire_599[ 6 ] = fresh_wire_714[ 6 ];
	assign fresh_wire_599[ 7 ] = fresh_wire_714[ 7 ];
	assign fresh_wire_599[ 8 ] = fresh_wire_714[ 8 ];
	assign fresh_wire_599[ 9 ] = fresh_wire_714[ 9 ];
	assign fresh_wire_599[ 10 ] = fresh_wire_714[ 10 ];
	assign fresh_wire_599[ 11 ] = fresh_wire_714[ 11 ];
	assign fresh_wire_599[ 12 ] = fresh_wire_714[ 12 ];
	assign fresh_wire_599[ 13 ] = fresh_wire_714[ 13 ];
	assign fresh_wire_599[ 14 ] = fresh_wire_714[ 14 ];
	assign fresh_wire_599[ 15 ] = fresh_wire_714[ 15 ];
	assign fresh_wire_599[ 16 ] = fresh_wire_714[ 16 ];
	assign fresh_wire_599[ 17 ] = fresh_wire_714[ 17 ];
	assign fresh_wire_599[ 18 ] = fresh_wire_714[ 18 ];
	assign fresh_wire_599[ 19 ] = fresh_wire_714[ 19 ];
	assign fresh_wire_599[ 20 ] = fresh_wire_714[ 20 ];
	assign fresh_wire_599[ 21 ] = fresh_wire_714[ 21 ];
	assign fresh_wire_599[ 22 ] = fresh_wire_714[ 22 ];
	assign fresh_wire_599[ 23 ] = fresh_wire_714[ 23 ];
	assign fresh_wire_599[ 24 ] = fresh_wire_714[ 24 ];
	assign fresh_wire_599[ 25 ] = fresh_wire_714[ 25 ];
	assign fresh_wire_599[ 26 ] = fresh_wire_714[ 26 ];
	assign fresh_wire_599[ 27 ] = fresh_wire_714[ 27 ];
	assign fresh_wire_599[ 28 ] = fresh_wire_714[ 28 ];
	assign fresh_wire_599[ 29 ] = fresh_wire_714[ 29 ];
	assign fresh_wire_599[ 30 ] = fresh_wire_714[ 30 ];
	assign fresh_wire_599[ 31 ] = fresh_wire_714[ 31 ];
	assign fresh_wire_601[ 0 ] = fresh_wire_216[ 0 ];
	assign fresh_wire_602[ 0 ] = fresh_wire_192[ 0 ];
	assign fresh_wire_602[ 1 ] = fresh_wire_192[ 1 ];
	assign fresh_wire_602[ 2 ] = fresh_wire_192[ 2 ];
	assign fresh_wire_602[ 3 ] = fresh_wire_192[ 3 ];
	assign fresh_wire_602[ 4 ] = fresh_wire_192[ 4 ];
	assign fresh_wire_602[ 5 ] = fresh_wire_192[ 5 ];
	assign fresh_wire_602[ 6 ] = fresh_wire_192[ 6 ];
	assign fresh_wire_602[ 7 ] = fresh_wire_192[ 7 ];
	assign fresh_wire_602[ 8 ] = fresh_wire_192[ 8 ];
	assign fresh_wire_602[ 9 ] = fresh_wire_192[ 9 ];
	assign fresh_wire_602[ 10 ] = fresh_wire_192[ 10 ];
	assign fresh_wire_602[ 11 ] = fresh_wire_192[ 11 ];
	assign fresh_wire_602[ 12 ] = fresh_wire_192[ 12 ];
	assign fresh_wire_602[ 13 ] = fresh_wire_192[ 13 ];
	assign fresh_wire_602[ 14 ] = fresh_wire_192[ 14 ];
	assign fresh_wire_602[ 15 ] = fresh_wire_192[ 15 ];
	assign fresh_wire_603[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_603[ 1 ] = fresh_wire_606[ 0 ];
	assign fresh_wire_603[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_603[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_603[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_603[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_603[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_603[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_603[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_603[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_603[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_603[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_603[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_603[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_603[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_603[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_605[ 0 ] = fresh_wire_243[ 0 ];
	assign fresh_wire_607[ 0 ] = fresh_wire_878[ 0 ];
	assign fresh_wire_607[ 1 ] = fresh_wire_878[ 1 ];
	assign fresh_wire_607[ 2 ] = fresh_wire_878[ 2 ];
	assign fresh_wire_607[ 3 ] = fresh_wire_878[ 3 ];
	assign fresh_wire_607[ 4 ] = fresh_wire_878[ 4 ];
	assign fresh_wire_607[ 5 ] = fresh_wire_878[ 5 ];
	assign fresh_wire_607[ 6 ] = fresh_wire_878[ 6 ];
	assign fresh_wire_607[ 7 ] = fresh_wire_878[ 7 ];
	assign fresh_wire_607[ 8 ] = fresh_wire_878[ 8 ];
	assign fresh_wire_607[ 9 ] = fresh_wire_878[ 9 ];
	assign fresh_wire_607[ 10 ] = fresh_wire_878[ 10 ];
	assign fresh_wire_607[ 11 ] = fresh_wire_878[ 11 ];
	assign fresh_wire_607[ 12 ] = fresh_wire_878[ 12 ];
	assign fresh_wire_607[ 13 ] = fresh_wire_878[ 13 ];
	assign fresh_wire_607[ 14 ] = fresh_wire_878[ 14 ];
	assign fresh_wire_607[ 15 ] = fresh_wire_878[ 15 ];
	assign fresh_wire_608[ 0 ] = fresh_wire_379[ 0 ];
	assign fresh_wire_608[ 1 ] = fresh_wire_379[ 1 ];
	assign fresh_wire_608[ 2 ] = fresh_wire_379[ 2 ];
	assign fresh_wire_608[ 3 ] = fresh_wire_379[ 3 ];
	assign fresh_wire_608[ 4 ] = fresh_wire_379[ 4 ];
	assign fresh_wire_608[ 5 ] = fresh_wire_379[ 5 ];
	assign fresh_wire_608[ 6 ] = fresh_wire_379[ 6 ];
	assign fresh_wire_608[ 7 ] = fresh_wire_379[ 7 ];
	assign fresh_wire_608[ 8 ] = fresh_wire_379[ 8 ];
	assign fresh_wire_608[ 9 ] = fresh_wire_379[ 9 ];
	assign fresh_wire_608[ 10 ] = fresh_wire_379[ 10 ];
	assign fresh_wire_608[ 11 ] = fresh_wire_379[ 11 ];
	assign fresh_wire_608[ 12 ] = fresh_wire_379[ 12 ];
	assign fresh_wire_608[ 13 ] = fresh_wire_379[ 13 ];
	assign fresh_wire_608[ 14 ] = fresh_wire_379[ 14 ];
	assign fresh_wire_608[ 15 ] = fresh_wire_379[ 15 ];
	assign fresh_wire_610[ 0 ] = fresh_wire_258[ 0 ];
	assign fresh_wire_611[ 0 ] = fresh_wire_666[ 0 ];
	assign fresh_wire_611[ 1 ] = fresh_wire_666[ 1 ];
	assign fresh_wire_612[ 0 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_612[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_614[ 0 ] = fresh_wire_426[ 0 ];
	assign fresh_wire_615[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_617[ 0 ] = fresh_wire_422[ 0 ];
	assign fresh_wire_618[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_620[ 0 ] = fresh_wire_426[ 0 ];
	assign fresh_wire_621[ 0 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_623[ 0 ] = fresh_wire_666[ 0 ];
	assign fresh_wire_623[ 1 ] = fresh_wire_666[ 1 ];
	assign fresh_wire_624[ 0 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_624[ 1 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_626[ 0 ] = fresh_wire_666[ 0 ];
	assign fresh_wire_626[ 1 ] = fresh_wire_666[ 1 ];
	assign fresh_wire_627[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_627[ 1 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_629[ 0 ] = fresh_wire_422[ 0 ];
	assign fresh_wire_630[ 0 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_632[ 0 ] = fresh_wire_666[ 0 ];
	assign fresh_wire_632[ 1 ] = fresh_wire_666[ 1 ];
	assign fresh_wire_633[ 0 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_633[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_635[ 0 ] = fresh_wire_666[ 0 ];
	assign fresh_wire_635[ 1 ] = fresh_wire_666[ 1 ];
	assign fresh_wire_636[ 0 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_636[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_638[ 0 ] = fresh_wire_616[ 0 ];
	assign fresh_wire_640[ 0 ] = fresh_wire_639[ 0 ];
	assign fresh_wire_641[ 0 ] = fresh_wire_644[ 0 ];
	assign fresh_wire_643[ 0 ] = fresh_wire_619[ 0 ];
	assign fresh_wire_645[ 0 ] = fresh_wire_2275[ 0 ];
	assign fresh_wire_646[ 0 ] = fresh_wire_649[ 0 ];
	assign fresh_wire_648[ 0 ] = fresh_wire_642[ 0 ];
	assign fresh_wire_650[ 0 ] = fresh_wire_2276[ 0 ];
	assign fresh_wire_651[ 0 ] = fresh_wire_654[ 0 ];
	assign fresh_wire_653[ 0 ] = fresh_wire_622[ 0 ];
	assign fresh_wire_655[ 0 ] = fresh_wire_2277[ 0 ];
	assign fresh_wire_656[ 0 ] = fresh_wire_659[ 0 ];
	assign fresh_wire_658[ 0 ] = fresh_wire_616[ 0 ];
	assign fresh_wire_660[ 0 ] = fresh_wire_2278[ 0 ];
	assign fresh_wire_661[ 0 ] = fresh_wire_664[ 0 ];
	assign fresh_wire_663[ 0 ] = fresh_wire_622[ 0 ];
	assign fresh_wire_665[ 0 ] = fresh_wire_686[ 0 ];
	assign fresh_wire_665[ 1 ] = fresh_wire_686[ 1 ];
	assign fresh_wire_667[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_668[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_669[ 0 ] = fresh_wire_96[ 0 ];
	assign fresh_wire_669[ 1 ] = fresh_wire_94[ 0 ];
	assign fresh_wire_669[ 2 ] = fresh_wire_92[ 0 ];
	assign fresh_wire_669[ 3 ] = fresh_wire_90[ 0 ];
	assign fresh_wire_669[ 4 ] = fresh_wire_88[ 0 ];
	assign fresh_wire_669[ 5 ] = fresh_wire_86[ 0 ];
	assign fresh_wire_669[ 6 ] = fresh_wire_114[ 0 ];
	assign fresh_wire_669[ 7 ] = fresh_wire_112[ 0 ];
	assign fresh_wire_669[ 8 ] = fresh_wire_110[ 0 ];
	assign fresh_wire_669[ 9 ] = fresh_wire_108[ 0 ];
	assign fresh_wire_669[ 10 ] = fresh_wire_106[ 0 ];
	assign fresh_wire_669[ 11 ] = fresh_wire_104[ 0 ];
	assign fresh_wire_669[ 12 ] = fresh_wire_102[ 0 ];
	assign fresh_wire_669[ 13 ] = fresh_wire_100[ 0 ];
	assign fresh_wire_669[ 14 ] = fresh_wire_98[ 0 ];
	assign fresh_wire_669[ 15 ] = fresh_wire_84[ 0 ];
	assign fresh_wire_669[ 16 ] = fresh_wire_670[ 0 ];
	assign fresh_wire_669[ 17 ] = fresh_wire_670[ 1 ];
	assign fresh_wire_669[ 18 ] = fresh_wire_670[ 2 ];
	assign fresh_wire_669[ 19 ] = fresh_wire_670[ 3 ];
	assign fresh_wire_669[ 20 ] = fresh_wire_670[ 4 ];
	assign fresh_wire_669[ 21 ] = fresh_wire_670[ 5 ];
	assign fresh_wire_669[ 22 ] = fresh_wire_670[ 6 ];
	assign fresh_wire_669[ 23 ] = fresh_wire_670[ 7 ];
	assign fresh_wire_669[ 24 ] = fresh_wire_670[ 8 ];
	assign fresh_wire_669[ 25 ] = fresh_wire_670[ 9 ];
	assign fresh_wire_669[ 26 ] = fresh_wire_670[ 10 ];
	assign fresh_wire_669[ 27 ] = fresh_wire_670[ 11 ];
	assign fresh_wire_669[ 28 ] = fresh_wire_670[ 12 ];
	assign fresh_wire_669[ 29 ] = fresh_wire_670[ 13 ];
	assign fresh_wire_669[ 30 ] = fresh_wire_670[ 14 ];
	assign fresh_wire_669[ 31 ] = fresh_wire_670[ 15 ];
	assign fresh_wire_669[ 32 ] = fresh_wire_670[ 16 ];
	assign fresh_wire_669[ 33 ] = fresh_wire_670[ 17 ];
	assign fresh_wire_669[ 34 ] = fresh_wire_670[ 18 ];
	assign fresh_wire_669[ 35 ] = fresh_wire_670[ 19 ];
	assign fresh_wire_669[ 36 ] = fresh_wire_670[ 20 ];
	assign fresh_wire_669[ 37 ] = fresh_wire_670[ 21 ];
	assign fresh_wire_669[ 38 ] = fresh_wire_670[ 22 ];
	assign fresh_wire_669[ 39 ] = fresh_wire_670[ 23 ];
	assign fresh_wire_669[ 40 ] = fresh_wire_670[ 24 ];
	assign fresh_wire_669[ 41 ] = fresh_wire_670[ 25 ];
	assign fresh_wire_669[ 42 ] = fresh_wire_670[ 26 ];
	assign fresh_wire_669[ 43 ] = fresh_wire_670[ 27 ];
	assign fresh_wire_669[ 44 ] = fresh_wire_670[ 28 ];
	assign fresh_wire_669[ 45 ] = fresh_wire_670[ 29 ];
	assign fresh_wire_669[ 46 ] = fresh_wire_670[ 30 ];
	assign fresh_wire_669[ 47 ] = fresh_wire_670[ 31 ];
	assign fresh_wire_671[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_672[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_673[ 0 ] = fresh_wire_625[ 0 ];
	assign fresh_wire_675[ 0 ] = fresh_wire_662[ 0 ];
	assign fresh_wire_676[ 0 ] = fresh_wire_674[ 0 ];
	assign fresh_wire_677[ 0 ] = fresh_wire_637[ 0 ];
	assign fresh_wire_679[ 0 ] = fresh_wire_657[ 0 ];
	assign fresh_wire_680[ 0 ] = fresh_wire_666[ 0 ];
	assign fresh_wire_680[ 1 ] = fresh_wire_666[ 1 ];
	assign fresh_wire_681[ 0 ] = fresh_wire_718[ 0 ];
	assign fresh_wire_681[ 1 ] = fresh_wire_718[ 1 ];
	assign fresh_wire_683[ 0 ] = fresh_wire_652[ 0 ];
	assign fresh_wire_684[ 0 ] = fresh_wire_682[ 0 ];
	assign fresh_wire_684[ 1 ] = fresh_wire_682[ 1 ];
	assign fresh_wire_685[ 0 ] = fresh_wire_613[ 0 ];
	assign fresh_wire_685[ 1 ] = fresh_wire_613[ 1 ];
	assign fresh_wire_687[ 0 ] = fresh_wire_647[ 0 ];
	assign fresh_wire_688[ 0 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 1 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 2 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 3 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 4 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 5 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 6 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 7 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 8 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 9 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 10 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 11 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 12 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 13 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 14 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 15 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 16 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 17 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 18 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 19 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 20 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 21 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 22 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 23 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 24 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 25 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 26 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 27 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 28 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 29 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 30 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_688[ 31 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_689[ 0 ] = fresh_wire_670[ 32 ];
	assign fresh_wire_689[ 1 ] = fresh_wire_670[ 33 ];
	assign fresh_wire_689[ 2 ] = fresh_wire_670[ 34 ];
	assign fresh_wire_689[ 3 ] = fresh_wire_670[ 35 ];
	assign fresh_wire_689[ 4 ] = fresh_wire_670[ 36 ];
	assign fresh_wire_689[ 5 ] = fresh_wire_670[ 37 ];
	assign fresh_wire_689[ 6 ] = fresh_wire_670[ 38 ];
	assign fresh_wire_689[ 7 ] = fresh_wire_670[ 39 ];
	assign fresh_wire_689[ 8 ] = fresh_wire_670[ 40 ];
	assign fresh_wire_689[ 9 ] = fresh_wire_670[ 41 ];
	assign fresh_wire_689[ 10 ] = fresh_wire_670[ 42 ];
	assign fresh_wire_689[ 11 ] = fresh_wire_670[ 43 ];
	assign fresh_wire_689[ 12 ] = fresh_wire_670[ 44 ];
	assign fresh_wire_689[ 13 ] = fresh_wire_670[ 45 ];
	assign fresh_wire_689[ 14 ] = fresh_wire_670[ 46 ];
	assign fresh_wire_689[ 15 ] = fresh_wire_670[ 47 ];
	assign fresh_wire_689[ 16 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_689[ 17 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_689[ 18 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_689[ 19 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_689[ 20 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_689[ 21 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_689[ 22 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_689[ 23 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_689[ 24 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_689[ 25 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_689[ 26 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_689[ 27 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_689[ 28 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_689[ 29 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_689[ 30 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_689[ 31 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_691[ 0 ] = fresh_wire_625[ 0 ];
	assign fresh_wire_692[ 0 ] = fresh_wire_690[ 0 ];
	assign fresh_wire_692[ 1 ] = fresh_wire_690[ 1 ];
	assign fresh_wire_692[ 2 ] = fresh_wire_690[ 2 ];
	assign fresh_wire_692[ 3 ] = fresh_wire_690[ 3 ];
	assign fresh_wire_692[ 4 ] = fresh_wire_690[ 4 ];
	assign fresh_wire_692[ 5 ] = fresh_wire_690[ 5 ];
	assign fresh_wire_692[ 6 ] = fresh_wire_690[ 6 ];
	assign fresh_wire_692[ 7 ] = fresh_wire_690[ 7 ];
	assign fresh_wire_692[ 8 ] = fresh_wire_690[ 8 ];
	assign fresh_wire_692[ 9 ] = fresh_wire_690[ 9 ];
	assign fresh_wire_692[ 10 ] = fresh_wire_690[ 10 ];
	assign fresh_wire_692[ 11 ] = fresh_wire_690[ 11 ];
	assign fresh_wire_692[ 12 ] = fresh_wire_690[ 12 ];
	assign fresh_wire_692[ 13 ] = fresh_wire_690[ 13 ];
	assign fresh_wire_692[ 14 ] = fresh_wire_690[ 14 ];
	assign fresh_wire_692[ 15 ] = fresh_wire_690[ 15 ];
	assign fresh_wire_692[ 16 ] = fresh_wire_690[ 16 ];
	assign fresh_wire_692[ 17 ] = fresh_wire_690[ 17 ];
	assign fresh_wire_692[ 18 ] = fresh_wire_690[ 18 ];
	assign fresh_wire_692[ 19 ] = fresh_wire_690[ 19 ];
	assign fresh_wire_692[ 20 ] = fresh_wire_690[ 20 ];
	assign fresh_wire_692[ 21 ] = fresh_wire_690[ 21 ];
	assign fresh_wire_692[ 22 ] = fresh_wire_690[ 22 ];
	assign fresh_wire_692[ 23 ] = fresh_wire_690[ 23 ];
	assign fresh_wire_692[ 24 ] = fresh_wire_690[ 24 ];
	assign fresh_wire_692[ 25 ] = fresh_wire_690[ 25 ];
	assign fresh_wire_692[ 26 ] = fresh_wire_690[ 26 ];
	assign fresh_wire_692[ 27 ] = fresh_wire_690[ 27 ];
	assign fresh_wire_692[ 28 ] = fresh_wire_690[ 28 ];
	assign fresh_wire_692[ 29 ] = fresh_wire_690[ 29 ];
	assign fresh_wire_692[ 30 ] = fresh_wire_690[ 30 ];
	assign fresh_wire_692[ 31 ] = fresh_wire_690[ 31 ];
	assign fresh_wire_693[ 0 ] = fresh_wire_670[ 16 ];
	assign fresh_wire_693[ 1 ] = fresh_wire_670[ 17 ];
	assign fresh_wire_693[ 2 ] = fresh_wire_670[ 18 ];
	assign fresh_wire_693[ 3 ] = fresh_wire_670[ 19 ];
	assign fresh_wire_693[ 4 ] = fresh_wire_670[ 20 ];
	assign fresh_wire_693[ 5 ] = fresh_wire_670[ 21 ];
	assign fresh_wire_693[ 6 ] = fresh_wire_670[ 22 ];
	assign fresh_wire_693[ 7 ] = fresh_wire_670[ 23 ];
	assign fresh_wire_693[ 8 ] = fresh_wire_670[ 24 ];
	assign fresh_wire_693[ 9 ] = fresh_wire_670[ 25 ];
	assign fresh_wire_693[ 10 ] = fresh_wire_670[ 26 ];
	assign fresh_wire_693[ 11 ] = fresh_wire_670[ 27 ];
	assign fresh_wire_693[ 12 ] = fresh_wire_670[ 28 ];
	assign fresh_wire_693[ 13 ] = fresh_wire_670[ 29 ];
	assign fresh_wire_693[ 14 ] = fresh_wire_670[ 30 ];
	assign fresh_wire_693[ 15 ] = fresh_wire_670[ 31 ];
	assign fresh_wire_693[ 16 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_693[ 17 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_693[ 18 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_693[ 19 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_693[ 20 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_693[ 21 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_693[ 22 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_693[ 23 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_693[ 24 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_693[ 25 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_693[ 26 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_693[ 27 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_693[ 28 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_693[ 29 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_693[ 30 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_693[ 31 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_695[ 0 ] = fresh_wire_628[ 0 ];
	assign fresh_wire_696[ 0 ] = fresh_wire_694[ 0 ];
	assign fresh_wire_696[ 1 ] = fresh_wire_694[ 1 ];
	assign fresh_wire_696[ 2 ] = fresh_wire_694[ 2 ];
	assign fresh_wire_696[ 3 ] = fresh_wire_694[ 3 ];
	assign fresh_wire_696[ 4 ] = fresh_wire_694[ 4 ];
	assign fresh_wire_696[ 5 ] = fresh_wire_694[ 5 ];
	assign fresh_wire_696[ 6 ] = fresh_wire_694[ 6 ];
	assign fresh_wire_696[ 7 ] = fresh_wire_694[ 7 ];
	assign fresh_wire_696[ 8 ] = fresh_wire_694[ 8 ];
	assign fresh_wire_696[ 9 ] = fresh_wire_694[ 9 ];
	assign fresh_wire_696[ 10 ] = fresh_wire_694[ 10 ];
	assign fresh_wire_696[ 11 ] = fresh_wire_694[ 11 ];
	assign fresh_wire_696[ 12 ] = fresh_wire_694[ 12 ];
	assign fresh_wire_696[ 13 ] = fresh_wire_694[ 13 ];
	assign fresh_wire_696[ 14 ] = fresh_wire_694[ 14 ];
	assign fresh_wire_696[ 15 ] = fresh_wire_694[ 15 ];
	assign fresh_wire_696[ 16 ] = fresh_wire_694[ 16 ];
	assign fresh_wire_696[ 17 ] = fresh_wire_694[ 17 ];
	assign fresh_wire_696[ 18 ] = fresh_wire_694[ 18 ];
	assign fresh_wire_696[ 19 ] = fresh_wire_694[ 19 ];
	assign fresh_wire_696[ 20 ] = fresh_wire_694[ 20 ];
	assign fresh_wire_696[ 21 ] = fresh_wire_694[ 21 ];
	assign fresh_wire_696[ 22 ] = fresh_wire_694[ 22 ];
	assign fresh_wire_696[ 23 ] = fresh_wire_694[ 23 ];
	assign fresh_wire_696[ 24 ] = fresh_wire_694[ 24 ];
	assign fresh_wire_696[ 25 ] = fresh_wire_694[ 25 ];
	assign fresh_wire_696[ 26 ] = fresh_wire_694[ 26 ];
	assign fresh_wire_696[ 27 ] = fresh_wire_694[ 27 ];
	assign fresh_wire_696[ 28 ] = fresh_wire_694[ 28 ];
	assign fresh_wire_696[ 29 ] = fresh_wire_694[ 29 ];
	assign fresh_wire_696[ 30 ] = fresh_wire_694[ 30 ];
	assign fresh_wire_696[ 31 ] = fresh_wire_694[ 31 ];
	assign fresh_wire_697[ 0 ] = fresh_wire_670[ 0 ];
	assign fresh_wire_697[ 1 ] = fresh_wire_670[ 1 ];
	assign fresh_wire_697[ 2 ] = fresh_wire_670[ 2 ];
	assign fresh_wire_697[ 3 ] = fresh_wire_670[ 3 ];
	assign fresh_wire_697[ 4 ] = fresh_wire_670[ 4 ];
	assign fresh_wire_697[ 5 ] = fresh_wire_670[ 5 ];
	assign fresh_wire_697[ 6 ] = fresh_wire_670[ 6 ];
	assign fresh_wire_697[ 7 ] = fresh_wire_670[ 7 ];
	assign fresh_wire_697[ 8 ] = fresh_wire_670[ 8 ];
	assign fresh_wire_697[ 9 ] = fresh_wire_670[ 9 ];
	assign fresh_wire_697[ 10 ] = fresh_wire_670[ 10 ];
	assign fresh_wire_697[ 11 ] = fresh_wire_670[ 11 ];
	assign fresh_wire_697[ 12 ] = fresh_wire_670[ 12 ];
	assign fresh_wire_697[ 13 ] = fresh_wire_670[ 13 ];
	assign fresh_wire_697[ 14 ] = fresh_wire_670[ 14 ];
	assign fresh_wire_697[ 15 ] = fresh_wire_670[ 15 ];
	assign fresh_wire_697[ 16 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_697[ 17 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_697[ 18 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_697[ 19 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_697[ 20 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_697[ 21 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_697[ 22 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_697[ 23 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_697[ 24 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_697[ 25 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_697[ 26 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_697[ 27 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_697[ 28 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_697[ 29 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_697[ 30 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_697[ 31 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_699[ 0 ] = fresh_wire_634[ 0 ];
	assign fresh_wire_700[ 0 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 1 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 2 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 3 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 4 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 5 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 6 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 7 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 8 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 9 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 10 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 11 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 12 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 13 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 14 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 15 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 16 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 17 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 18 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 19 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 20 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 21 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 22 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 23 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 24 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 25 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 26 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 27 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 28 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 29 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 30 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_700[ 31 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_701[ 0 ] = fresh_wire_698[ 0 ];
	assign fresh_wire_701[ 1 ] = fresh_wire_698[ 1 ];
	assign fresh_wire_701[ 2 ] = fresh_wire_698[ 2 ];
	assign fresh_wire_701[ 3 ] = fresh_wire_698[ 3 ];
	assign fresh_wire_701[ 4 ] = fresh_wire_698[ 4 ];
	assign fresh_wire_701[ 5 ] = fresh_wire_698[ 5 ];
	assign fresh_wire_701[ 6 ] = fresh_wire_698[ 6 ];
	assign fresh_wire_701[ 7 ] = fresh_wire_698[ 7 ];
	assign fresh_wire_701[ 8 ] = fresh_wire_698[ 8 ];
	assign fresh_wire_701[ 9 ] = fresh_wire_698[ 9 ];
	assign fresh_wire_701[ 10 ] = fresh_wire_698[ 10 ];
	assign fresh_wire_701[ 11 ] = fresh_wire_698[ 11 ];
	assign fresh_wire_701[ 12 ] = fresh_wire_698[ 12 ];
	assign fresh_wire_701[ 13 ] = fresh_wire_698[ 13 ];
	assign fresh_wire_701[ 14 ] = fresh_wire_698[ 14 ];
	assign fresh_wire_701[ 15 ] = fresh_wire_698[ 15 ];
	assign fresh_wire_701[ 16 ] = fresh_wire_698[ 16 ];
	assign fresh_wire_701[ 17 ] = fresh_wire_698[ 17 ];
	assign fresh_wire_701[ 18 ] = fresh_wire_698[ 18 ];
	assign fresh_wire_701[ 19 ] = fresh_wire_698[ 19 ];
	assign fresh_wire_701[ 20 ] = fresh_wire_698[ 20 ];
	assign fresh_wire_701[ 21 ] = fresh_wire_698[ 21 ];
	assign fresh_wire_701[ 22 ] = fresh_wire_698[ 22 ];
	assign fresh_wire_701[ 23 ] = fresh_wire_698[ 23 ];
	assign fresh_wire_701[ 24 ] = fresh_wire_698[ 24 ];
	assign fresh_wire_701[ 25 ] = fresh_wire_698[ 25 ];
	assign fresh_wire_701[ 26 ] = fresh_wire_698[ 26 ];
	assign fresh_wire_701[ 27 ] = fresh_wire_698[ 27 ];
	assign fresh_wire_701[ 28 ] = fresh_wire_698[ 28 ];
	assign fresh_wire_701[ 29 ] = fresh_wire_698[ 29 ];
	assign fresh_wire_701[ 30 ] = fresh_wire_698[ 30 ];
	assign fresh_wire_701[ 31 ] = fresh_wire_698[ 31 ];
	assign fresh_wire_703[ 0 ] = fresh_wire_631[ 0 ];
	assign fresh_wire_704[ 0 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 1 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 2 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 3 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 4 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 5 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 6 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 7 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 8 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 9 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 10 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 11 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 12 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 13 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 14 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 15 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 16 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 17 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 18 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 19 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 20 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 21 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 22 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 23 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 24 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 25 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 26 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 27 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 28 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 29 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 30 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_704[ 31 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_705[ 0 ] = fresh_wire_670[ 16 ];
	assign fresh_wire_705[ 1 ] = fresh_wire_670[ 17 ];
	assign fresh_wire_705[ 2 ] = fresh_wire_670[ 18 ];
	assign fresh_wire_705[ 3 ] = fresh_wire_670[ 19 ];
	assign fresh_wire_705[ 4 ] = fresh_wire_670[ 20 ];
	assign fresh_wire_705[ 5 ] = fresh_wire_670[ 21 ];
	assign fresh_wire_705[ 6 ] = fresh_wire_670[ 22 ];
	assign fresh_wire_705[ 7 ] = fresh_wire_670[ 23 ];
	assign fresh_wire_705[ 8 ] = fresh_wire_670[ 24 ];
	assign fresh_wire_705[ 9 ] = fresh_wire_670[ 25 ];
	assign fresh_wire_705[ 10 ] = fresh_wire_670[ 26 ];
	assign fresh_wire_705[ 11 ] = fresh_wire_670[ 27 ];
	assign fresh_wire_705[ 12 ] = fresh_wire_670[ 28 ];
	assign fresh_wire_705[ 13 ] = fresh_wire_670[ 29 ];
	assign fresh_wire_705[ 14 ] = fresh_wire_670[ 30 ];
	assign fresh_wire_705[ 15 ] = fresh_wire_670[ 31 ];
	assign fresh_wire_705[ 16 ] = fresh_wire_670[ 32 ];
	assign fresh_wire_705[ 17 ] = fresh_wire_670[ 33 ];
	assign fresh_wire_705[ 18 ] = fresh_wire_670[ 34 ];
	assign fresh_wire_705[ 19 ] = fresh_wire_670[ 35 ];
	assign fresh_wire_705[ 20 ] = fresh_wire_670[ 36 ];
	assign fresh_wire_705[ 21 ] = fresh_wire_670[ 37 ];
	assign fresh_wire_705[ 22 ] = fresh_wire_670[ 38 ];
	assign fresh_wire_705[ 23 ] = fresh_wire_670[ 39 ];
	assign fresh_wire_705[ 24 ] = fresh_wire_670[ 40 ];
	assign fresh_wire_705[ 25 ] = fresh_wire_670[ 41 ];
	assign fresh_wire_705[ 26 ] = fresh_wire_670[ 42 ];
	assign fresh_wire_705[ 27 ] = fresh_wire_670[ 43 ];
	assign fresh_wire_705[ 28 ] = fresh_wire_670[ 44 ];
	assign fresh_wire_705[ 29 ] = fresh_wire_670[ 45 ];
	assign fresh_wire_705[ 30 ] = fresh_wire_670[ 46 ];
	assign fresh_wire_705[ 31 ] = fresh_wire_670[ 47 ];
	assign fresh_wire_707[ 0 ] = fresh_wire_625[ 0 ];
	assign fresh_wire_708[ 0 ] = fresh_wire_706[ 0 ];
	assign fresh_wire_708[ 1 ] = fresh_wire_706[ 1 ];
	assign fresh_wire_708[ 2 ] = fresh_wire_706[ 2 ];
	assign fresh_wire_708[ 3 ] = fresh_wire_706[ 3 ];
	assign fresh_wire_708[ 4 ] = fresh_wire_706[ 4 ];
	assign fresh_wire_708[ 5 ] = fresh_wire_706[ 5 ];
	assign fresh_wire_708[ 6 ] = fresh_wire_706[ 6 ];
	assign fresh_wire_708[ 7 ] = fresh_wire_706[ 7 ];
	assign fresh_wire_708[ 8 ] = fresh_wire_706[ 8 ];
	assign fresh_wire_708[ 9 ] = fresh_wire_706[ 9 ];
	assign fresh_wire_708[ 10 ] = fresh_wire_706[ 10 ];
	assign fresh_wire_708[ 11 ] = fresh_wire_706[ 11 ];
	assign fresh_wire_708[ 12 ] = fresh_wire_706[ 12 ];
	assign fresh_wire_708[ 13 ] = fresh_wire_706[ 13 ];
	assign fresh_wire_708[ 14 ] = fresh_wire_706[ 14 ];
	assign fresh_wire_708[ 15 ] = fresh_wire_706[ 15 ];
	assign fresh_wire_708[ 16 ] = fresh_wire_706[ 16 ];
	assign fresh_wire_708[ 17 ] = fresh_wire_706[ 17 ];
	assign fresh_wire_708[ 18 ] = fresh_wire_706[ 18 ];
	assign fresh_wire_708[ 19 ] = fresh_wire_706[ 19 ];
	assign fresh_wire_708[ 20 ] = fresh_wire_706[ 20 ];
	assign fresh_wire_708[ 21 ] = fresh_wire_706[ 21 ];
	assign fresh_wire_708[ 22 ] = fresh_wire_706[ 22 ];
	assign fresh_wire_708[ 23 ] = fresh_wire_706[ 23 ];
	assign fresh_wire_708[ 24 ] = fresh_wire_706[ 24 ];
	assign fresh_wire_708[ 25 ] = fresh_wire_706[ 25 ];
	assign fresh_wire_708[ 26 ] = fresh_wire_706[ 26 ];
	assign fresh_wire_708[ 27 ] = fresh_wire_706[ 27 ];
	assign fresh_wire_708[ 28 ] = fresh_wire_706[ 28 ];
	assign fresh_wire_708[ 29 ] = fresh_wire_706[ 29 ];
	assign fresh_wire_708[ 30 ] = fresh_wire_706[ 30 ];
	assign fresh_wire_708[ 31 ] = fresh_wire_706[ 31 ];
	assign fresh_wire_709[ 0 ] = fresh_wire_670[ 0 ];
	assign fresh_wire_709[ 1 ] = fresh_wire_670[ 1 ];
	assign fresh_wire_709[ 2 ] = fresh_wire_670[ 2 ];
	assign fresh_wire_709[ 3 ] = fresh_wire_670[ 3 ];
	assign fresh_wire_709[ 4 ] = fresh_wire_670[ 4 ];
	assign fresh_wire_709[ 5 ] = fresh_wire_670[ 5 ];
	assign fresh_wire_709[ 6 ] = fresh_wire_670[ 6 ];
	assign fresh_wire_709[ 7 ] = fresh_wire_670[ 7 ];
	assign fresh_wire_709[ 8 ] = fresh_wire_670[ 8 ];
	assign fresh_wire_709[ 9 ] = fresh_wire_670[ 9 ];
	assign fresh_wire_709[ 10 ] = fresh_wire_670[ 10 ];
	assign fresh_wire_709[ 11 ] = fresh_wire_670[ 11 ];
	assign fresh_wire_709[ 12 ] = fresh_wire_670[ 12 ];
	assign fresh_wire_709[ 13 ] = fresh_wire_670[ 13 ];
	assign fresh_wire_709[ 14 ] = fresh_wire_670[ 14 ];
	assign fresh_wire_709[ 15 ] = fresh_wire_670[ 15 ];
	assign fresh_wire_709[ 16 ] = fresh_wire_670[ 16 ];
	assign fresh_wire_709[ 17 ] = fresh_wire_670[ 17 ];
	assign fresh_wire_709[ 18 ] = fresh_wire_670[ 18 ];
	assign fresh_wire_709[ 19 ] = fresh_wire_670[ 19 ];
	assign fresh_wire_709[ 20 ] = fresh_wire_670[ 20 ];
	assign fresh_wire_709[ 21 ] = fresh_wire_670[ 21 ];
	assign fresh_wire_709[ 22 ] = fresh_wire_670[ 22 ];
	assign fresh_wire_709[ 23 ] = fresh_wire_670[ 23 ];
	assign fresh_wire_709[ 24 ] = fresh_wire_670[ 24 ];
	assign fresh_wire_709[ 25 ] = fresh_wire_670[ 25 ];
	assign fresh_wire_709[ 26 ] = fresh_wire_670[ 26 ];
	assign fresh_wire_709[ 27 ] = fresh_wire_670[ 27 ];
	assign fresh_wire_709[ 28 ] = fresh_wire_670[ 28 ];
	assign fresh_wire_709[ 29 ] = fresh_wire_670[ 29 ];
	assign fresh_wire_709[ 30 ] = fresh_wire_670[ 30 ];
	assign fresh_wire_709[ 31 ] = fresh_wire_670[ 31 ];
	assign fresh_wire_711[ 0 ] = fresh_wire_628[ 0 ];
	assign fresh_wire_712[ 0 ] = fresh_wire_702[ 0 ];
	assign fresh_wire_712[ 1 ] = fresh_wire_702[ 1 ];
	assign fresh_wire_712[ 2 ] = fresh_wire_702[ 2 ];
	assign fresh_wire_712[ 3 ] = fresh_wire_702[ 3 ];
	assign fresh_wire_712[ 4 ] = fresh_wire_702[ 4 ];
	assign fresh_wire_712[ 5 ] = fresh_wire_702[ 5 ];
	assign fresh_wire_712[ 6 ] = fresh_wire_702[ 6 ];
	assign fresh_wire_712[ 7 ] = fresh_wire_702[ 7 ];
	assign fresh_wire_712[ 8 ] = fresh_wire_702[ 8 ];
	assign fresh_wire_712[ 9 ] = fresh_wire_702[ 9 ];
	assign fresh_wire_712[ 10 ] = fresh_wire_702[ 10 ];
	assign fresh_wire_712[ 11 ] = fresh_wire_702[ 11 ];
	assign fresh_wire_712[ 12 ] = fresh_wire_702[ 12 ];
	assign fresh_wire_712[ 13 ] = fresh_wire_702[ 13 ];
	assign fresh_wire_712[ 14 ] = fresh_wire_702[ 14 ];
	assign fresh_wire_712[ 15 ] = fresh_wire_702[ 15 ];
	assign fresh_wire_712[ 16 ] = fresh_wire_702[ 16 ];
	assign fresh_wire_712[ 17 ] = fresh_wire_702[ 17 ];
	assign fresh_wire_712[ 18 ] = fresh_wire_702[ 18 ];
	assign fresh_wire_712[ 19 ] = fresh_wire_702[ 19 ];
	assign fresh_wire_712[ 20 ] = fresh_wire_702[ 20 ];
	assign fresh_wire_712[ 21 ] = fresh_wire_702[ 21 ];
	assign fresh_wire_712[ 22 ] = fresh_wire_702[ 22 ];
	assign fresh_wire_712[ 23 ] = fresh_wire_702[ 23 ];
	assign fresh_wire_712[ 24 ] = fresh_wire_702[ 24 ];
	assign fresh_wire_712[ 25 ] = fresh_wire_702[ 25 ];
	assign fresh_wire_712[ 26 ] = fresh_wire_702[ 26 ];
	assign fresh_wire_712[ 27 ] = fresh_wire_702[ 27 ];
	assign fresh_wire_712[ 28 ] = fresh_wire_702[ 28 ];
	assign fresh_wire_712[ 29 ] = fresh_wire_702[ 29 ];
	assign fresh_wire_712[ 30 ] = fresh_wire_702[ 30 ];
	assign fresh_wire_712[ 31 ] = fresh_wire_702[ 31 ];
	assign fresh_wire_713[ 0 ] = fresh_wire_710[ 0 ];
	assign fresh_wire_713[ 1 ] = fresh_wire_710[ 1 ];
	assign fresh_wire_713[ 2 ] = fresh_wire_710[ 2 ];
	assign fresh_wire_713[ 3 ] = fresh_wire_710[ 3 ];
	assign fresh_wire_713[ 4 ] = fresh_wire_710[ 4 ];
	assign fresh_wire_713[ 5 ] = fresh_wire_710[ 5 ];
	assign fresh_wire_713[ 6 ] = fresh_wire_710[ 6 ];
	assign fresh_wire_713[ 7 ] = fresh_wire_710[ 7 ];
	assign fresh_wire_713[ 8 ] = fresh_wire_710[ 8 ];
	assign fresh_wire_713[ 9 ] = fresh_wire_710[ 9 ];
	assign fresh_wire_713[ 10 ] = fresh_wire_710[ 10 ];
	assign fresh_wire_713[ 11 ] = fresh_wire_710[ 11 ];
	assign fresh_wire_713[ 12 ] = fresh_wire_710[ 12 ];
	assign fresh_wire_713[ 13 ] = fresh_wire_710[ 13 ];
	assign fresh_wire_713[ 14 ] = fresh_wire_710[ 14 ];
	assign fresh_wire_713[ 15 ] = fresh_wire_710[ 15 ];
	assign fresh_wire_713[ 16 ] = fresh_wire_710[ 16 ];
	assign fresh_wire_713[ 17 ] = fresh_wire_710[ 17 ];
	assign fresh_wire_713[ 18 ] = fresh_wire_710[ 18 ];
	assign fresh_wire_713[ 19 ] = fresh_wire_710[ 19 ];
	assign fresh_wire_713[ 20 ] = fresh_wire_710[ 20 ];
	assign fresh_wire_713[ 21 ] = fresh_wire_710[ 21 ];
	assign fresh_wire_713[ 22 ] = fresh_wire_710[ 22 ];
	assign fresh_wire_713[ 23 ] = fresh_wire_710[ 23 ];
	assign fresh_wire_713[ 24 ] = fresh_wire_710[ 24 ];
	assign fresh_wire_713[ 25 ] = fresh_wire_710[ 25 ];
	assign fresh_wire_713[ 26 ] = fresh_wire_710[ 26 ];
	assign fresh_wire_713[ 27 ] = fresh_wire_710[ 27 ];
	assign fresh_wire_713[ 28 ] = fresh_wire_710[ 28 ];
	assign fresh_wire_713[ 29 ] = fresh_wire_710[ 29 ];
	assign fresh_wire_713[ 30 ] = fresh_wire_710[ 30 ];
	assign fresh_wire_713[ 31 ] = fresh_wire_710[ 31 ];
	assign fresh_wire_715[ 0 ] = fresh_wire_622[ 0 ];
	assign fresh_wire_716[ 0 ] = fresh_wire_666[ 0 ];
	assign fresh_wire_716[ 1 ] = fresh_wire_666[ 1 ];
	assign fresh_wire_717[ 0 ] = fresh_wire_719[ 0 ];
	assign fresh_wire_717[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_720[ 0 ] = fresh_wire_858[ 0 ];
	assign fresh_wire_720[ 1 ] = fresh_wire_858[ 1 ];
	assign fresh_wire_721[ 0 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_721[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_723[ 0 ] = fresh_wire_858[ 0 ];
	assign fresh_wire_723[ 1 ] = fresh_wire_858[ 1 ];
	assign fresh_wire_724[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_724[ 1 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_726[ 0 ] = fresh_wire_386[ 0 ];
	assign fresh_wire_727[ 0 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_729[ 0 ] = fresh_wire_382[ 0 ];
	assign fresh_wire_730[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_732[ 0 ] = fresh_wire_390[ 0 ];
	assign fresh_wire_733[ 0 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_735[ 0 ] = fresh_wire_382[ 0 ];
	assign fresh_wire_736[ 0 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_738[ 0 ] = fresh_wire_386[ 0 ];
	assign fresh_wire_739[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_741[ 0 ] = fresh_wire_390[ 0 ];
	assign fresh_wire_742[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_744[ 0 ] = fresh_wire_858[ 0 ];
	assign fresh_wire_744[ 1 ] = fresh_wire_858[ 1 ];
	assign fresh_wire_745[ 0 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_745[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_747[ 0 ] = fresh_wire_858[ 0 ];
	assign fresh_wire_747[ 1 ] = fresh_wire_858[ 1 ];
	assign fresh_wire_748[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_748[ 1 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_750[ 0 ] = fresh_wire_858[ 0 ];
	assign fresh_wire_750[ 1 ] = fresh_wire_858[ 1 ];
	assign fresh_wire_751[ 0 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_751[ 1 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_753[ 0 ] = fresh_wire_858[ 0 ];
	assign fresh_wire_753[ 1 ] = fresh_wire_858[ 1 ];
	assign fresh_wire_754[ 0 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_754[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_756[ 0 ] = fresh_wire_858[ 0 ];
	assign fresh_wire_756[ 1 ] = fresh_wire_858[ 1 ];
	assign fresh_wire_757[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_757[ 1 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_759[ 0 ] = fresh_wire_728[ 0 ];
	assign fresh_wire_761[ 0 ] = fresh_wire_760[ 0 ];
	assign fresh_wire_762[ 0 ] = fresh_wire_765[ 0 ];
	assign fresh_wire_764[ 0 ] = fresh_wire_731[ 0 ];
	assign fresh_wire_766[ 0 ] = fresh_wire_734[ 0 ];
	assign fresh_wire_768[ 0 ] = fresh_wire_767[ 0 ];
	assign fresh_wire_769[ 0 ] = fresh_wire_772[ 0 ];
	assign fresh_wire_771[ 0 ] = fresh_wire_731[ 0 ];
	assign fresh_wire_773[ 0 ] = fresh_wire_728[ 0 ];
	assign fresh_wire_775[ 0 ] = fresh_wire_774[ 0 ];
	assign fresh_wire_776[ 0 ] = fresh_wire_779[ 0 ];
	assign fresh_wire_778[ 0 ] = fresh_wire_737[ 0 ];
	assign fresh_wire_780[ 0 ] = fresh_wire_734[ 0 ];
	assign fresh_wire_782[ 0 ] = fresh_wire_781[ 0 ];
	assign fresh_wire_783[ 0 ] = fresh_wire_786[ 0 ];
	assign fresh_wire_785[ 0 ] = fresh_wire_737[ 0 ];
	assign fresh_wire_787[ 0 ] = fresh_wire_740[ 0 ];
	assign fresh_wire_789[ 0 ] = fresh_wire_788[ 0 ];
	assign fresh_wire_790[ 0 ] = fresh_wire_793[ 0 ];
	assign fresh_wire_792[ 0 ] = fresh_wire_743[ 0 ];
	assign fresh_wire_794[ 0 ] = fresh_wire_791[ 0 ];
	assign fresh_wire_796[ 0 ] = fresh_wire_795[ 0 ];
	assign fresh_wire_797[ 0 ] = fresh_wire_800[ 0 ];
	assign fresh_wire_799[ 0 ] = fresh_wire_731[ 0 ];
	assign fresh_wire_801[ 0 ] = fresh_wire_740[ 0 ];
	assign fresh_wire_803[ 0 ] = fresh_wire_802[ 0 ];
	assign fresh_wire_804[ 0 ] = fresh_wire_807[ 0 ];
	assign fresh_wire_806[ 0 ] = fresh_wire_743[ 0 ];
	assign fresh_wire_808[ 0 ] = fresh_wire_805[ 0 ];
	assign fresh_wire_810[ 0 ] = fresh_wire_809[ 0 ];
	assign fresh_wire_811[ 0 ] = fresh_wire_814[ 0 ];
	assign fresh_wire_813[ 0 ] = fresh_wire_737[ 0 ];
	assign fresh_wire_815[ 0 ] = fresh_wire_849[ 0 ];
	assign fresh_wire_817[ 0 ] = fresh_wire_816[ 0 ];
	assign fresh_wire_818[ 0 ] = fresh_wire_821[ 0 ];
	assign fresh_wire_820[ 0 ] = fresh_wire_731[ 0 ];
	assign fresh_wire_822[ 0 ] = fresh_wire_856[ 0 ];
	assign fresh_wire_824[ 0 ] = fresh_wire_823[ 0 ];
	assign fresh_wire_825[ 0 ] = fresh_wire_828[ 0 ];
	assign fresh_wire_827[ 0 ] = fresh_wire_737[ 0 ];
	assign fresh_wire_829[ 0 ] = fresh_wire_740[ 0 ];
	assign fresh_wire_831[ 0 ] = fresh_wire_830[ 0 ];
	assign fresh_wire_832[ 0 ] = fresh_wire_835[ 0 ];
	assign fresh_wire_834[ 0 ] = fresh_wire_743[ 0 ];
	assign fresh_wire_836[ 0 ] = fresh_wire_833[ 0 ];
	assign fresh_wire_838[ 0 ] = fresh_wire_837[ 0 ];
	assign fresh_wire_839[ 0 ] = fresh_wire_842[ 0 ];
	assign fresh_wire_841[ 0 ] = fresh_wire_737[ 0 ];
	assign fresh_wire_843[ 0 ] = fresh_wire_728[ 0 ];
	assign fresh_wire_845[ 0 ] = fresh_wire_734[ 0 ];
	assign fresh_wire_847[ 0 ] = fresh_wire_844[ 0 ];
	assign fresh_wire_848[ 0 ] = fresh_wire_846[ 0 ];
	assign fresh_wire_850[ 0 ] = fresh_wire_728[ 0 ];
	assign fresh_wire_852[ 0 ] = fresh_wire_734[ 0 ];
	assign fresh_wire_854[ 0 ] = fresh_wire_851[ 0 ];
	assign fresh_wire_855[ 0 ] = fresh_wire_853[ 0 ];
	assign fresh_wire_857[ 0 ] = fresh_wire_914[ 0 ];
	assign fresh_wire_857[ 1 ] = fresh_wire_914[ 1 ];
	assign fresh_wire_859[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_860[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_861[ 0 ] = fresh_wire_922[ 0 ];
	assign fresh_wire_861[ 1 ] = fresh_wire_922[ 1 ];
	assign fresh_wire_861[ 2 ] = fresh_wire_922[ 2 ];
	assign fresh_wire_861[ 3 ] = fresh_wire_922[ 3 ];
	assign fresh_wire_861[ 4 ] = fresh_wire_922[ 4 ];
	assign fresh_wire_861[ 5 ] = fresh_wire_922[ 5 ];
	assign fresh_wire_861[ 6 ] = fresh_wire_922[ 6 ];
	assign fresh_wire_861[ 7 ] = fresh_wire_922[ 7 ];
	assign fresh_wire_861[ 8 ] = fresh_wire_922[ 8 ];
	assign fresh_wire_861[ 9 ] = fresh_wire_922[ 9 ];
	assign fresh_wire_861[ 10 ] = fresh_wire_922[ 10 ];
	assign fresh_wire_861[ 11 ] = fresh_wire_922[ 11 ];
	assign fresh_wire_861[ 12 ] = fresh_wire_922[ 12 ];
	assign fresh_wire_861[ 13 ] = fresh_wire_922[ 13 ];
	assign fresh_wire_861[ 14 ] = fresh_wire_922[ 14 ];
	assign fresh_wire_861[ 15 ] = fresh_wire_922[ 15 ];
	assign fresh_wire_861[ 16 ] = fresh_wire_922[ 16 ];
	assign fresh_wire_861[ 17 ] = fresh_wire_922[ 17 ];
	assign fresh_wire_861[ 18 ] = fresh_wire_922[ 18 ];
	assign fresh_wire_861[ 19 ] = fresh_wire_922[ 19 ];
	assign fresh_wire_861[ 20 ] = fresh_wire_922[ 20 ];
	assign fresh_wire_861[ 21 ] = fresh_wire_922[ 21 ];
	assign fresh_wire_861[ 22 ] = fresh_wire_922[ 22 ];
	assign fresh_wire_861[ 23 ] = fresh_wire_922[ 23 ];
	assign fresh_wire_861[ 24 ] = fresh_wire_922[ 24 ];
	assign fresh_wire_861[ 25 ] = fresh_wire_922[ 25 ];
	assign fresh_wire_861[ 26 ] = fresh_wire_922[ 26 ];
	assign fresh_wire_861[ 27 ] = fresh_wire_922[ 27 ];
	assign fresh_wire_861[ 28 ] = fresh_wire_922[ 28 ];
	assign fresh_wire_861[ 29 ] = fresh_wire_922[ 29 ];
	assign fresh_wire_861[ 30 ] = fresh_wire_922[ 30 ];
	assign fresh_wire_861[ 31 ] = fresh_wire_922[ 31 ];
	assign fresh_wire_861[ 32 ] = fresh_wire_922[ 32 ];
	assign fresh_wire_861[ 33 ] = fresh_wire_922[ 33 ];
	assign fresh_wire_861[ 34 ] = fresh_wire_922[ 34 ];
	assign fresh_wire_861[ 35 ] = fresh_wire_922[ 35 ];
	assign fresh_wire_861[ 36 ] = fresh_wire_922[ 36 ];
	assign fresh_wire_861[ 37 ] = fresh_wire_922[ 37 ];
	assign fresh_wire_861[ 38 ] = fresh_wire_922[ 38 ];
	assign fresh_wire_861[ 39 ] = fresh_wire_922[ 39 ];
	assign fresh_wire_861[ 40 ] = fresh_wire_922[ 40 ];
	assign fresh_wire_861[ 41 ] = fresh_wire_922[ 41 ];
	assign fresh_wire_861[ 42 ] = fresh_wire_922[ 42 ];
	assign fresh_wire_861[ 43 ] = fresh_wire_922[ 43 ];
	assign fresh_wire_861[ 44 ] = fresh_wire_922[ 44 ];
	assign fresh_wire_861[ 45 ] = fresh_wire_922[ 45 ];
	assign fresh_wire_861[ 46 ] = fresh_wire_922[ 46 ];
	assign fresh_wire_861[ 47 ] = fresh_wire_922[ 47 ];
	assign fresh_wire_863[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_864[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_864[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_864[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_864[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_864[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_864[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_864[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_864[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_864[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_864[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_864[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_864[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_864[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_864[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_864[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_864[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_865[ 0 ] = fresh_wire_862[ 32 ];
	assign fresh_wire_865[ 1 ] = fresh_wire_862[ 33 ];
	assign fresh_wire_865[ 2 ] = fresh_wire_862[ 34 ];
	assign fresh_wire_865[ 3 ] = fresh_wire_862[ 35 ];
	assign fresh_wire_865[ 4 ] = fresh_wire_862[ 36 ];
	assign fresh_wire_865[ 5 ] = fresh_wire_862[ 37 ];
	assign fresh_wire_865[ 6 ] = fresh_wire_862[ 38 ];
	assign fresh_wire_865[ 7 ] = fresh_wire_862[ 39 ];
	assign fresh_wire_865[ 8 ] = fresh_wire_862[ 40 ];
	assign fresh_wire_865[ 9 ] = fresh_wire_862[ 41 ];
	assign fresh_wire_865[ 10 ] = fresh_wire_862[ 42 ];
	assign fresh_wire_865[ 11 ] = fresh_wire_862[ 43 ];
	assign fresh_wire_865[ 12 ] = fresh_wire_862[ 44 ];
	assign fresh_wire_865[ 13 ] = fresh_wire_862[ 45 ];
	assign fresh_wire_865[ 14 ] = fresh_wire_862[ 46 ];
	assign fresh_wire_865[ 15 ] = fresh_wire_862[ 47 ];
	assign fresh_wire_867[ 0 ] = fresh_wire_752[ 0 ];
	assign fresh_wire_868[ 0 ] = fresh_wire_866[ 0 ];
	assign fresh_wire_868[ 1 ] = fresh_wire_866[ 1 ];
	assign fresh_wire_868[ 2 ] = fresh_wire_866[ 2 ];
	assign fresh_wire_868[ 3 ] = fresh_wire_866[ 3 ];
	assign fresh_wire_868[ 4 ] = fresh_wire_866[ 4 ];
	assign fresh_wire_868[ 5 ] = fresh_wire_866[ 5 ];
	assign fresh_wire_868[ 6 ] = fresh_wire_866[ 6 ];
	assign fresh_wire_868[ 7 ] = fresh_wire_866[ 7 ];
	assign fresh_wire_868[ 8 ] = fresh_wire_866[ 8 ];
	assign fresh_wire_868[ 9 ] = fresh_wire_866[ 9 ];
	assign fresh_wire_868[ 10 ] = fresh_wire_866[ 10 ];
	assign fresh_wire_868[ 11 ] = fresh_wire_866[ 11 ];
	assign fresh_wire_868[ 12 ] = fresh_wire_866[ 12 ];
	assign fresh_wire_868[ 13 ] = fresh_wire_866[ 13 ];
	assign fresh_wire_868[ 14 ] = fresh_wire_866[ 14 ];
	assign fresh_wire_868[ 15 ] = fresh_wire_866[ 15 ];
	assign fresh_wire_869[ 0 ] = fresh_wire_862[ 16 ];
	assign fresh_wire_869[ 1 ] = fresh_wire_862[ 17 ];
	assign fresh_wire_869[ 2 ] = fresh_wire_862[ 18 ];
	assign fresh_wire_869[ 3 ] = fresh_wire_862[ 19 ];
	assign fresh_wire_869[ 4 ] = fresh_wire_862[ 20 ];
	assign fresh_wire_869[ 5 ] = fresh_wire_862[ 21 ];
	assign fresh_wire_869[ 6 ] = fresh_wire_862[ 22 ];
	assign fresh_wire_869[ 7 ] = fresh_wire_862[ 23 ];
	assign fresh_wire_869[ 8 ] = fresh_wire_862[ 24 ];
	assign fresh_wire_869[ 9 ] = fresh_wire_862[ 25 ];
	assign fresh_wire_869[ 10 ] = fresh_wire_862[ 26 ];
	assign fresh_wire_869[ 11 ] = fresh_wire_862[ 27 ];
	assign fresh_wire_869[ 12 ] = fresh_wire_862[ 28 ];
	assign fresh_wire_869[ 13 ] = fresh_wire_862[ 29 ];
	assign fresh_wire_869[ 14 ] = fresh_wire_862[ 30 ];
	assign fresh_wire_869[ 15 ] = fresh_wire_862[ 31 ];
	assign fresh_wire_871[ 0 ] = fresh_wire_749[ 0 ];
	assign fresh_wire_872[ 0 ] = fresh_wire_870[ 0 ];
	assign fresh_wire_872[ 1 ] = fresh_wire_870[ 1 ];
	assign fresh_wire_872[ 2 ] = fresh_wire_870[ 2 ];
	assign fresh_wire_872[ 3 ] = fresh_wire_870[ 3 ];
	assign fresh_wire_872[ 4 ] = fresh_wire_870[ 4 ];
	assign fresh_wire_872[ 5 ] = fresh_wire_870[ 5 ];
	assign fresh_wire_872[ 6 ] = fresh_wire_870[ 6 ];
	assign fresh_wire_872[ 7 ] = fresh_wire_870[ 7 ];
	assign fresh_wire_872[ 8 ] = fresh_wire_870[ 8 ];
	assign fresh_wire_872[ 9 ] = fresh_wire_870[ 9 ];
	assign fresh_wire_872[ 10 ] = fresh_wire_870[ 10 ];
	assign fresh_wire_872[ 11 ] = fresh_wire_870[ 11 ];
	assign fresh_wire_872[ 12 ] = fresh_wire_870[ 12 ];
	assign fresh_wire_872[ 13 ] = fresh_wire_870[ 13 ];
	assign fresh_wire_872[ 14 ] = fresh_wire_870[ 14 ];
	assign fresh_wire_872[ 15 ] = fresh_wire_870[ 15 ];
	assign fresh_wire_873[ 0 ] = fresh_wire_862[ 0 ];
	assign fresh_wire_873[ 1 ] = fresh_wire_862[ 1 ];
	assign fresh_wire_873[ 2 ] = fresh_wire_862[ 2 ];
	assign fresh_wire_873[ 3 ] = fresh_wire_862[ 3 ];
	assign fresh_wire_873[ 4 ] = fresh_wire_862[ 4 ];
	assign fresh_wire_873[ 5 ] = fresh_wire_862[ 5 ];
	assign fresh_wire_873[ 6 ] = fresh_wire_862[ 6 ];
	assign fresh_wire_873[ 7 ] = fresh_wire_862[ 7 ];
	assign fresh_wire_873[ 8 ] = fresh_wire_862[ 8 ];
	assign fresh_wire_873[ 9 ] = fresh_wire_862[ 9 ];
	assign fresh_wire_873[ 10 ] = fresh_wire_862[ 10 ];
	assign fresh_wire_873[ 11 ] = fresh_wire_862[ 11 ];
	assign fresh_wire_873[ 12 ] = fresh_wire_862[ 12 ];
	assign fresh_wire_873[ 13 ] = fresh_wire_862[ 13 ];
	assign fresh_wire_873[ 14 ] = fresh_wire_862[ 14 ];
	assign fresh_wire_873[ 15 ] = fresh_wire_862[ 15 ];
	assign fresh_wire_875[ 0 ] = fresh_wire_746[ 0 ];
	assign fresh_wire_876[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_876[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_876[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_876[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_876[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_876[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_876[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_876[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_876[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_876[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_876[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_876[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_876[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_876[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_876[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_876[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_877[ 0 ] = fresh_wire_874[ 0 ];
	assign fresh_wire_877[ 1 ] = fresh_wire_874[ 1 ];
	assign fresh_wire_877[ 2 ] = fresh_wire_874[ 2 ];
	assign fresh_wire_877[ 3 ] = fresh_wire_874[ 3 ];
	assign fresh_wire_877[ 4 ] = fresh_wire_874[ 4 ];
	assign fresh_wire_877[ 5 ] = fresh_wire_874[ 5 ];
	assign fresh_wire_877[ 6 ] = fresh_wire_874[ 6 ];
	assign fresh_wire_877[ 7 ] = fresh_wire_874[ 7 ];
	assign fresh_wire_877[ 8 ] = fresh_wire_874[ 8 ];
	assign fresh_wire_877[ 9 ] = fresh_wire_874[ 9 ];
	assign fresh_wire_877[ 10 ] = fresh_wire_874[ 10 ];
	assign fresh_wire_877[ 11 ] = fresh_wire_874[ 11 ];
	assign fresh_wire_877[ 12 ] = fresh_wire_874[ 12 ];
	assign fresh_wire_877[ 13 ] = fresh_wire_874[ 13 ];
	assign fresh_wire_877[ 14 ] = fresh_wire_874[ 14 ];
	assign fresh_wire_877[ 15 ] = fresh_wire_874[ 15 ];
	assign fresh_wire_879[ 0 ] = fresh_wire_737[ 0 ];
	assign fresh_wire_880[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_881[ 0 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_883[ 0 ] = fresh_wire_826[ 0 ];
	assign fresh_wire_884[ 0 ] = fresh_wire_882[ 0 ];
	assign fresh_wire_885[ 0 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_887[ 0 ] = fresh_wire_819[ 0 ];
	assign fresh_wire_888[ 0 ] = fresh_wire_886[ 0 ];
	assign fresh_wire_889[ 0 ] = fresh_wire_758[ 0 ];
	assign fresh_wire_891[ 0 ] = fresh_wire_812[ 0 ];
	assign fresh_wire_892[ 0 ] = fresh_wire_890[ 0 ];
	assign fresh_wire_893[ 0 ] = fresh_wire_755[ 0 ];
	assign fresh_wire_895[ 0 ] = fresh_wire_798[ 0 ];
	assign fresh_wire_896[ 0 ] = fresh_wire_858[ 0 ];
	assign fresh_wire_896[ 1 ] = fresh_wire_858[ 1 ];
	assign fresh_wire_897[ 0 ] = fresh_wire_722[ 0 ];
	assign fresh_wire_897[ 1 ] = fresh_wire_722[ 1 ];
	assign fresh_wire_899[ 0 ] = fresh_wire_784[ 0 ];
	assign fresh_wire_900[ 0 ] = fresh_wire_898[ 0 ];
	assign fresh_wire_900[ 1 ] = fresh_wire_898[ 1 ];
	assign fresh_wire_901[ 0 ] = fresh_wire_858[ 0 ];
	assign fresh_wire_901[ 1 ] = fresh_wire_858[ 1 ];
	assign fresh_wire_903[ 0 ] = fresh_wire_777[ 0 ];
	assign fresh_wire_904[ 0 ] = fresh_wire_902[ 0 ];
	assign fresh_wire_904[ 1 ] = fresh_wire_902[ 1 ];
	assign fresh_wire_905[ 0 ] = fresh_wire_725[ 0 ];
	assign fresh_wire_905[ 1 ] = fresh_wire_725[ 1 ];
	assign fresh_wire_907[ 0 ] = fresh_wire_770[ 0 ];
	assign fresh_wire_908[ 0 ] = fresh_wire_906[ 0 ];
	assign fresh_wire_908[ 1 ] = fresh_wire_906[ 1 ];
	assign fresh_wire_909[ 0 ] = fresh_wire_722[ 0 ];
	assign fresh_wire_909[ 1 ] = fresh_wire_722[ 1 ];
	assign fresh_wire_911[ 0 ] = fresh_wire_763[ 0 ];
	assign fresh_wire_912[ 0 ] = fresh_wire_910[ 0 ];
	assign fresh_wire_912[ 1 ] = fresh_wire_910[ 1 ];
	assign fresh_wire_913[ 0 ] = fresh_wire_926[ 0 ];
	assign fresh_wire_913[ 1 ] = fresh_wire_926[ 1 ];
	assign fresh_wire_915[ 0 ] = fresh_wire_840[ 0 ];
	assign fresh_wire_916[ 0 ] = fresh_wire_862[ 0 ];
	assign fresh_wire_916[ 1 ] = fresh_wire_862[ 1 ];
	assign fresh_wire_916[ 2 ] = fresh_wire_862[ 2 ];
	assign fresh_wire_916[ 3 ] = fresh_wire_862[ 3 ];
	assign fresh_wire_916[ 4 ] = fresh_wire_862[ 4 ];
	assign fresh_wire_916[ 5 ] = fresh_wire_862[ 5 ];
	assign fresh_wire_916[ 6 ] = fresh_wire_862[ 6 ];
	assign fresh_wire_916[ 7 ] = fresh_wire_862[ 7 ];
	assign fresh_wire_916[ 8 ] = fresh_wire_862[ 8 ];
	assign fresh_wire_916[ 9 ] = fresh_wire_862[ 9 ];
	assign fresh_wire_916[ 10 ] = fresh_wire_862[ 10 ];
	assign fresh_wire_916[ 11 ] = fresh_wire_862[ 11 ];
	assign fresh_wire_916[ 12 ] = fresh_wire_862[ 12 ];
	assign fresh_wire_916[ 13 ] = fresh_wire_862[ 13 ];
	assign fresh_wire_916[ 14 ] = fresh_wire_862[ 14 ];
	assign fresh_wire_916[ 15 ] = fresh_wire_862[ 15 ];
	assign fresh_wire_916[ 16 ] = fresh_wire_862[ 16 ];
	assign fresh_wire_916[ 17 ] = fresh_wire_862[ 17 ];
	assign fresh_wire_916[ 18 ] = fresh_wire_862[ 18 ];
	assign fresh_wire_916[ 19 ] = fresh_wire_862[ 19 ];
	assign fresh_wire_916[ 20 ] = fresh_wire_862[ 20 ];
	assign fresh_wire_916[ 21 ] = fresh_wire_862[ 21 ];
	assign fresh_wire_916[ 22 ] = fresh_wire_862[ 22 ];
	assign fresh_wire_916[ 23 ] = fresh_wire_862[ 23 ];
	assign fresh_wire_916[ 24 ] = fresh_wire_862[ 24 ];
	assign fresh_wire_916[ 25 ] = fresh_wire_862[ 25 ];
	assign fresh_wire_916[ 26 ] = fresh_wire_862[ 26 ];
	assign fresh_wire_916[ 27 ] = fresh_wire_862[ 27 ];
	assign fresh_wire_916[ 28 ] = fresh_wire_862[ 28 ];
	assign fresh_wire_916[ 29 ] = fresh_wire_862[ 29 ];
	assign fresh_wire_916[ 30 ] = fresh_wire_862[ 30 ];
	assign fresh_wire_916[ 31 ] = fresh_wire_862[ 31 ];
	assign fresh_wire_916[ 32 ] = fresh_wire_862[ 32 ];
	assign fresh_wire_916[ 33 ] = fresh_wire_862[ 33 ];
	assign fresh_wire_916[ 34 ] = fresh_wire_862[ 34 ];
	assign fresh_wire_916[ 35 ] = fresh_wire_862[ 35 ];
	assign fresh_wire_916[ 36 ] = fresh_wire_862[ 36 ];
	assign fresh_wire_916[ 37 ] = fresh_wire_862[ 37 ];
	assign fresh_wire_916[ 38 ] = fresh_wire_862[ 38 ];
	assign fresh_wire_916[ 39 ] = fresh_wire_862[ 39 ];
	assign fresh_wire_916[ 40 ] = fresh_wire_862[ 40 ];
	assign fresh_wire_916[ 41 ] = fresh_wire_862[ 41 ];
	assign fresh_wire_916[ 42 ] = fresh_wire_862[ 42 ];
	assign fresh_wire_916[ 43 ] = fresh_wire_862[ 43 ];
	assign fresh_wire_916[ 44 ] = fresh_wire_862[ 44 ];
	assign fresh_wire_916[ 45 ] = fresh_wire_862[ 45 ];
	assign fresh_wire_916[ 46 ] = fresh_wire_862[ 46 ];
	assign fresh_wire_916[ 47 ] = fresh_wire_862[ 47 ];
	assign fresh_wire_917[ 0 ] = fresh_wire_600[ 0 ];
	assign fresh_wire_917[ 1 ] = fresh_wire_600[ 1 ];
	assign fresh_wire_917[ 2 ] = fresh_wire_600[ 2 ];
	assign fresh_wire_917[ 3 ] = fresh_wire_600[ 3 ];
	assign fresh_wire_917[ 4 ] = fresh_wire_600[ 4 ];
	assign fresh_wire_917[ 5 ] = fresh_wire_600[ 5 ];
	assign fresh_wire_917[ 6 ] = fresh_wire_600[ 6 ];
	assign fresh_wire_917[ 7 ] = fresh_wire_600[ 7 ];
	assign fresh_wire_917[ 8 ] = fresh_wire_600[ 8 ];
	assign fresh_wire_917[ 9 ] = fresh_wire_600[ 9 ];
	assign fresh_wire_917[ 10 ] = fresh_wire_600[ 10 ];
	assign fresh_wire_917[ 11 ] = fresh_wire_600[ 11 ];
	assign fresh_wire_917[ 12 ] = fresh_wire_600[ 12 ];
	assign fresh_wire_917[ 13 ] = fresh_wire_600[ 13 ];
	assign fresh_wire_917[ 14 ] = fresh_wire_600[ 14 ];
	assign fresh_wire_917[ 15 ] = fresh_wire_600[ 15 ];
	assign fresh_wire_917[ 16 ] = fresh_wire_862[ 0 ];
	assign fresh_wire_917[ 17 ] = fresh_wire_862[ 1 ];
	assign fresh_wire_917[ 18 ] = fresh_wire_862[ 2 ];
	assign fresh_wire_917[ 19 ] = fresh_wire_862[ 3 ];
	assign fresh_wire_917[ 20 ] = fresh_wire_862[ 4 ];
	assign fresh_wire_917[ 21 ] = fresh_wire_862[ 5 ];
	assign fresh_wire_917[ 22 ] = fresh_wire_862[ 6 ];
	assign fresh_wire_917[ 23 ] = fresh_wire_862[ 7 ];
	assign fresh_wire_917[ 24 ] = fresh_wire_862[ 8 ];
	assign fresh_wire_917[ 25 ] = fresh_wire_862[ 9 ];
	assign fresh_wire_917[ 26 ] = fresh_wire_862[ 10 ];
	assign fresh_wire_917[ 27 ] = fresh_wire_862[ 11 ];
	assign fresh_wire_917[ 28 ] = fresh_wire_862[ 12 ];
	assign fresh_wire_917[ 29 ] = fresh_wire_862[ 13 ];
	assign fresh_wire_917[ 30 ] = fresh_wire_862[ 14 ];
	assign fresh_wire_917[ 31 ] = fresh_wire_862[ 15 ];
	assign fresh_wire_917[ 32 ] = fresh_wire_862[ 16 ];
	assign fresh_wire_917[ 33 ] = fresh_wire_862[ 17 ];
	assign fresh_wire_917[ 34 ] = fresh_wire_862[ 18 ];
	assign fresh_wire_917[ 35 ] = fresh_wire_862[ 19 ];
	assign fresh_wire_917[ 36 ] = fresh_wire_862[ 20 ];
	assign fresh_wire_917[ 37 ] = fresh_wire_862[ 21 ];
	assign fresh_wire_917[ 38 ] = fresh_wire_862[ 22 ];
	assign fresh_wire_917[ 39 ] = fresh_wire_862[ 23 ];
	assign fresh_wire_917[ 40 ] = fresh_wire_862[ 24 ];
	assign fresh_wire_917[ 41 ] = fresh_wire_862[ 25 ];
	assign fresh_wire_917[ 42 ] = fresh_wire_862[ 26 ];
	assign fresh_wire_917[ 43 ] = fresh_wire_862[ 27 ];
	assign fresh_wire_917[ 44 ] = fresh_wire_862[ 28 ];
	assign fresh_wire_917[ 45 ] = fresh_wire_862[ 29 ];
	assign fresh_wire_917[ 46 ] = fresh_wire_862[ 30 ];
	assign fresh_wire_917[ 47 ] = fresh_wire_862[ 31 ];
	assign fresh_wire_919[ 0 ] = fresh_wire_728[ 0 ];
	assign fresh_wire_920[ 0 ] = fresh_wire_918[ 0 ];
	assign fresh_wire_920[ 1 ] = fresh_wire_918[ 1 ];
	assign fresh_wire_920[ 2 ] = fresh_wire_918[ 2 ];
	assign fresh_wire_920[ 3 ] = fresh_wire_918[ 3 ];
	assign fresh_wire_920[ 4 ] = fresh_wire_918[ 4 ];
	assign fresh_wire_920[ 5 ] = fresh_wire_918[ 5 ];
	assign fresh_wire_920[ 6 ] = fresh_wire_918[ 6 ];
	assign fresh_wire_920[ 7 ] = fresh_wire_918[ 7 ];
	assign fresh_wire_920[ 8 ] = fresh_wire_918[ 8 ];
	assign fresh_wire_920[ 9 ] = fresh_wire_918[ 9 ];
	assign fresh_wire_920[ 10 ] = fresh_wire_918[ 10 ];
	assign fresh_wire_920[ 11 ] = fresh_wire_918[ 11 ];
	assign fresh_wire_920[ 12 ] = fresh_wire_918[ 12 ];
	assign fresh_wire_920[ 13 ] = fresh_wire_918[ 13 ];
	assign fresh_wire_920[ 14 ] = fresh_wire_918[ 14 ];
	assign fresh_wire_920[ 15 ] = fresh_wire_918[ 15 ];
	assign fresh_wire_920[ 16 ] = fresh_wire_918[ 16 ];
	assign fresh_wire_920[ 17 ] = fresh_wire_918[ 17 ];
	assign fresh_wire_920[ 18 ] = fresh_wire_918[ 18 ];
	assign fresh_wire_920[ 19 ] = fresh_wire_918[ 19 ];
	assign fresh_wire_920[ 20 ] = fresh_wire_918[ 20 ];
	assign fresh_wire_920[ 21 ] = fresh_wire_918[ 21 ];
	assign fresh_wire_920[ 22 ] = fresh_wire_918[ 22 ];
	assign fresh_wire_920[ 23 ] = fresh_wire_918[ 23 ];
	assign fresh_wire_920[ 24 ] = fresh_wire_918[ 24 ];
	assign fresh_wire_920[ 25 ] = fresh_wire_918[ 25 ];
	assign fresh_wire_920[ 26 ] = fresh_wire_918[ 26 ];
	assign fresh_wire_920[ 27 ] = fresh_wire_918[ 27 ];
	assign fresh_wire_920[ 28 ] = fresh_wire_918[ 28 ];
	assign fresh_wire_920[ 29 ] = fresh_wire_918[ 29 ];
	assign fresh_wire_920[ 30 ] = fresh_wire_918[ 30 ];
	assign fresh_wire_920[ 31 ] = fresh_wire_918[ 31 ];
	assign fresh_wire_920[ 32 ] = fresh_wire_918[ 32 ];
	assign fresh_wire_920[ 33 ] = fresh_wire_918[ 33 ];
	assign fresh_wire_920[ 34 ] = fresh_wire_918[ 34 ];
	assign fresh_wire_920[ 35 ] = fresh_wire_918[ 35 ];
	assign fresh_wire_920[ 36 ] = fresh_wire_918[ 36 ];
	assign fresh_wire_920[ 37 ] = fresh_wire_918[ 37 ];
	assign fresh_wire_920[ 38 ] = fresh_wire_918[ 38 ];
	assign fresh_wire_920[ 39 ] = fresh_wire_918[ 39 ];
	assign fresh_wire_920[ 40 ] = fresh_wire_918[ 40 ];
	assign fresh_wire_920[ 41 ] = fresh_wire_918[ 41 ];
	assign fresh_wire_920[ 42 ] = fresh_wire_918[ 42 ];
	assign fresh_wire_920[ 43 ] = fresh_wire_918[ 43 ];
	assign fresh_wire_920[ 44 ] = fresh_wire_918[ 44 ];
	assign fresh_wire_920[ 45 ] = fresh_wire_918[ 45 ];
	assign fresh_wire_920[ 46 ] = fresh_wire_918[ 46 ];
	assign fresh_wire_920[ 47 ] = fresh_wire_918[ 47 ];
	assign fresh_wire_921[ 0 ] = fresh_wire_600[ 0 ];
	assign fresh_wire_921[ 1 ] = fresh_wire_600[ 1 ];
	assign fresh_wire_921[ 2 ] = fresh_wire_600[ 2 ];
	assign fresh_wire_921[ 3 ] = fresh_wire_600[ 3 ];
	assign fresh_wire_921[ 4 ] = fresh_wire_600[ 4 ];
	assign fresh_wire_921[ 5 ] = fresh_wire_600[ 5 ];
	assign fresh_wire_921[ 6 ] = fresh_wire_600[ 6 ];
	assign fresh_wire_921[ 7 ] = fresh_wire_600[ 7 ];
	assign fresh_wire_921[ 8 ] = fresh_wire_600[ 8 ];
	assign fresh_wire_921[ 9 ] = fresh_wire_600[ 9 ];
	assign fresh_wire_921[ 10 ] = fresh_wire_600[ 10 ];
	assign fresh_wire_921[ 11 ] = fresh_wire_600[ 11 ];
	assign fresh_wire_921[ 12 ] = fresh_wire_600[ 12 ];
	assign fresh_wire_921[ 13 ] = fresh_wire_600[ 13 ];
	assign fresh_wire_921[ 14 ] = fresh_wire_600[ 14 ];
	assign fresh_wire_921[ 15 ] = fresh_wire_600[ 15 ];
	assign fresh_wire_921[ 16 ] = fresh_wire_600[ 16 ];
	assign fresh_wire_921[ 17 ] = fresh_wire_600[ 17 ];
	assign fresh_wire_921[ 18 ] = fresh_wire_600[ 18 ];
	assign fresh_wire_921[ 19 ] = fresh_wire_600[ 19 ];
	assign fresh_wire_921[ 20 ] = fresh_wire_600[ 20 ];
	assign fresh_wire_921[ 21 ] = fresh_wire_600[ 21 ];
	assign fresh_wire_921[ 22 ] = fresh_wire_600[ 22 ];
	assign fresh_wire_921[ 23 ] = fresh_wire_600[ 23 ];
	assign fresh_wire_921[ 24 ] = fresh_wire_600[ 24 ];
	assign fresh_wire_921[ 25 ] = fresh_wire_600[ 25 ];
	assign fresh_wire_921[ 26 ] = fresh_wire_600[ 26 ];
	assign fresh_wire_921[ 27 ] = fresh_wire_600[ 27 ];
	assign fresh_wire_921[ 28 ] = fresh_wire_600[ 28 ];
	assign fresh_wire_921[ 29 ] = fresh_wire_600[ 29 ];
	assign fresh_wire_921[ 30 ] = fresh_wire_600[ 30 ];
	assign fresh_wire_921[ 31 ] = fresh_wire_600[ 31 ];
	assign fresh_wire_921[ 32 ] = fresh_wire_862[ 0 ];
	assign fresh_wire_921[ 33 ] = fresh_wire_862[ 1 ];
	assign fresh_wire_921[ 34 ] = fresh_wire_862[ 2 ];
	assign fresh_wire_921[ 35 ] = fresh_wire_862[ 3 ];
	assign fresh_wire_921[ 36 ] = fresh_wire_862[ 4 ];
	assign fresh_wire_921[ 37 ] = fresh_wire_862[ 5 ];
	assign fresh_wire_921[ 38 ] = fresh_wire_862[ 6 ];
	assign fresh_wire_921[ 39 ] = fresh_wire_862[ 7 ];
	assign fresh_wire_921[ 40 ] = fresh_wire_862[ 8 ];
	assign fresh_wire_921[ 41 ] = fresh_wire_862[ 9 ];
	assign fresh_wire_921[ 42 ] = fresh_wire_862[ 10 ];
	assign fresh_wire_921[ 43 ] = fresh_wire_862[ 11 ];
	assign fresh_wire_921[ 44 ] = fresh_wire_862[ 12 ];
	assign fresh_wire_921[ 45 ] = fresh_wire_862[ 13 ];
	assign fresh_wire_921[ 46 ] = fresh_wire_862[ 14 ];
	assign fresh_wire_921[ 47 ] = fresh_wire_862[ 15 ];
	assign fresh_wire_923[ 0 ] = fresh_wire_734[ 0 ];
	assign fresh_wire_924[ 0 ] = fresh_wire_858[ 0 ];
	assign fresh_wire_924[ 1 ] = fresh_wire_858[ 1 ];
	assign fresh_wire_925[ 0 ] = fresh_wire_927[ 0 ];
	assign fresh_wire_925[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_928[ 0 ] = fresh_wire_157[ 0 ];
	assign fresh_wire_930[ 0 ] = fresh_wire_426[ 0 ];
	assign fresh_wire_932[ 0 ] = fresh_wire_929[ 0 ];
	assign fresh_wire_933[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_935[ 0 ] = fresh_wire_931[ 0 ];
	assign fresh_wire_936[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_938[ 0 ] = fresh_wire_943[ 0 ];
	assign fresh_wire_938[ 1 ] = fresh_wire_943[ 1 ];
	assign fresh_wire_938[ 2 ] = fresh_wire_943[ 2 ];
	assign fresh_wire_938[ 3 ] = fresh_wire_943[ 3 ];
	assign fresh_wire_938[ 4 ] = fresh_wire_943[ 4 ];
	assign fresh_wire_938[ 5 ] = fresh_wire_943[ 5 ];
	assign fresh_wire_938[ 6 ] = fresh_wire_943[ 6 ];
	assign fresh_wire_938[ 7 ] = fresh_wire_943[ 7 ];
	assign fresh_wire_938[ 8 ] = fresh_wire_943[ 8 ];
	assign fresh_wire_938[ 9 ] = fresh_wire_943[ 9 ];
	assign fresh_wire_938[ 10 ] = fresh_wire_943[ 10 ];
	assign fresh_wire_938[ 11 ] = fresh_wire_943[ 11 ];
	assign fresh_wire_938[ 12 ] = fresh_wire_943[ 12 ];
	assign fresh_wire_938[ 13 ] = fresh_wire_943[ 13 ];
	assign fresh_wire_938[ 14 ] = fresh_wire_943[ 14 ];
	assign fresh_wire_938[ 15 ] = fresh_wire_943[ 15 ];
	assign fresh_wire_940[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_941[ 0 ] = fresh_wire_939[ 0 ];
	assign fresh_wire_941[ 1 ] = fresh_wire_939[ 1 ];
	assign fresh_wire_941[ 2 ] = fresh_wire_939[ 2 ];
	assign fresh_wire_941[ 3 ] = fresh_wire_939[ 3 ];
	assign fresh_wire_941[ 4 ] = fresh_wire_939[ 4 ];
	assign fresh_wire_941[ 5 ] = fresh_wire_939[ 5 ];
	assign fresh_wire_941[ 6 ] = fresh_wire_939[ 6 ];
	assign fresh_wire_941[ 7 ] = fresh_wire_939[ 7 ];
	assign fresh_wire_941[ 8 ] = fresh_wire_939[ 8 ];
	assign fresh_wire_941[ 9 ] = fresh_wire_939[ 9 ];
	assign fresh_wire_941[ 10 ] = fresh_wire_939[ 10 ];
	assign fresh_wire_941[ 11 ] = fresh_wire_939[ 11 ];
	assign fresh_wire_941[ 12 ] = fresh_wire_939[ 12 ];
	assign fresh_wire_941[ 13 ] = fresh_wire_939[ 13 ];
	assign fresh_wire_941[ 14 ] = fresh_wire_939[ 14 ];
	assign fresh_wire_941[ 15 ] = fresh_wire_939[ 15 ];
	assign fresh_wire_942[ 0 ] = fresh_wire_1022[ 0 ];
	assign fresh_wire_942[ 1 ] = fresh_wire_1022[ 1 ];
	assign fresh_wire_942[ 2 ] = fresh_wire_1022[ 2 ];
	assign fresh_wire_942[ 3 ] = fresh_wire_1022[ 3 ];
	assign fresh_wire_942[ 4 ] = fresh_wire_1022[ 4 ];
	assign fresh_wire_942[ 5 ] = fresh_wire_1022[ 5 ];
	assign fresh_wire_942[ 6 ] = fresh_wire_1022[ 6 ];
	assign fresh_wire_942[ 7 ] = fresh_wire_1022[ 7 ];
	assign fresh_wire_942[ 8 ] = fresh_wire_1022[ 8 ];
	assign fresh_wire_942[ 9 ] = fresh_wire_1022[ 9 ];
	assign fresh_wire_942[ 10 ] = fresh_wire_1022[ 10 ];
	assign fresh_wire_942[ 11 ] = fresh_wire_1022[ 11 ];
	assign fresh_wire_942[ 12 ] = fresh_wire_1022[ 12 ];
	assign fresh_wire_942[ 13 ] = fresh_wire_1022[ 13 ];
	assign fresh_wire_942[ 14 ] = fresh_wire_1022[ 14 ];
	assign fresh_wire_942[ 15 ] = fresh_wire_1022[ 15 ];
	assign fresh_wire_944[ 0 ] = fresh_wire_934[ 0 ];
	assign fresh_wire_945[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_945[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_945[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_945[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_945[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_945[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_945[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_945[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_945[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_945[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_945[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_945[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_945[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_945[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_945[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_945[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_946[ 0 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 1 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 2 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 3 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 4 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 5 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 6 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 7 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 8 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 9 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 10 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 11 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 12 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 13 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 14 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_946[ 15 ] = fresh_wire_949[ 0 ];
	assign fresh_wire_948[ 0 ] = fresh_wire_937[ 0 ];
	assign fresh_wire_950[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_950[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_950[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_950[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_950[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_950[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_950[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_950[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_950[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_950[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_950[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_950[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_950[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_950[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_950[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_950[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_951[ 0 ] = fresh_wire_947[ 0 ];
	assign fresh_wire_951[ 1 ] = fresh_wire_947[ 1 ];
	assign fresh_wire_951[ 2 ] = fresh_wire_947[ 2 ];
	assign fresh_wire_951[ 3 ] = fresh_wire_947[ 3 ];
	assign fresh_wire_951[ 4 ] = fresh_wire_947[ 4 ];
	assign fresh_wire_951[ 5 ] = fresh_wire_947[ 5 ];
	assign fresh_wire_951[ 6 ] = fresh_wire_947[ 6 ];
	assign fresh_wire_951[ 7 ] = fresh_wire_947[ 7 ];
	assign fresh_wire_951[ 8 ] = fresh_wire_947[ 8 ];
	assign fresh_wire_951[ 9 ] = fresh_wire_947[ 9 ];
	assign fresh_wire_951[ 10 ] = fresh_wire_947[ 10 ];
	assign fresh_wire_951[ 11 ] = fresh_wire_947[ 11 ];
	assign fresh_wire_951[ 12 ] = fresh_wire_947[ 12 ];
	assign fresh_wire_951[ 13 ] = fresh_wire_947[ 13 ];
	assign fresh_wire_951[ 14 ] = fresh_wire_947[ 14 ];
	assign fresh_wire_951[ 15 ] = fresh_wire_947[ 15 ];
	assign fresh_wire_953[ 0 ] = fresh_wire_934[ 0 ];
	assign fresh_wire_954[ 0 ] = fresh_wire_958[ 0 ];
	assign fresh_wire_954[ 1 ] = fresh_wire_965[ 0 ];
	assign fresh_wire_954[ 2 ] = fresh_wire_966[ 0 ];
	assign fresh_wire_954[ 3 ] = fresh_wire_967[ 0 ];
	assign fresh_wire_954[ 4 ] = fresh_wire_968[ 0 ];
	assign fresh_wire_954[ 5 ] = fresh_wire_969[ 0 ];
	assign fresh_wire_954[ 6 ] = fresh_wire_970[ 0 ];
	assign fresh_wire_954[ 7 ] = fresh_wire_971[ 0 ];
	assign fresh_wire_954[ 8 ] = fresh_wire_972[ 0 ];
	assign fresh_wire_954[ 9 ] = fresh_wire_973[ 0 ];
	assign fresh_wire_954[ 10 ] = fresh_wire_959[ 0 ];
	assign fresh_wire_954[ 11 ] = fresh_wire_960[ 0 ];
	assign fresh_wire_954[ 12 ] = fresh_wire_961[ 0 ];
	assign fresh_wire_954[ 13 ] = fresh_wire_962[ 0 ];
	assign fresh_wire_954[ 14 ] = fresh_wire_963[ 0 ];
	assign fresh_wire_954[ 15 ] = fresh_wire_964[ 0 ];
	assign fresh_wire_955[ 0 ] = fresh_wire_714[ 0 ];
	assign fresh_wire_955[ 1 ] = fresh_wire_714[ 1 ];
	assign fresh_wire_955[ 2 ] = fresh_wire_714[ 2 ];
	assign fresh_wire_955[ 3 ] = fresh_wire_714[ 3 ];
	assign fresh_wire_955[ 4 ] = fresh_wire_714[ 4 ];
	assign fresh_wire_955[ 5 ] = fresh_wire_714[ 5 ];
	assign fresh_wire_955[ 6 ] = fresh_wire_714[ 6 ];
	assign fresh_wire_955[ 7 ] = fresh_wire_714[ 7 ];
	assign fresh_wire_955[ 8 ] = fresh_wire_714[ 8 ];
	assign fresh_wire_955[ 9 ] = fresh_wire_714[ 9 ];
	assign fresh_wire_955[ 10 ] = fresh_wire_714[ 10 ];
	assign fresh_wire_955[ 11 ] = fresh_wire_714[ 11 ];
	assign fresh_wire_955[ 12 ] = fresh_wire_714[ 12 ];
	assign fresh_wire_955[ 13 ] = fresh_wire_714[ 13 ];
	assign fresh_wire_955[ 14 ] = fresh_wire_714[ 14 ];
	assign fresh_wire_955[ 15 ] = fresh_wire_714[ 15 ];
	assign fresh_wire_957[ 0 ] = fresh_wire_937[ 0 ];
	assign fresh_wire_974[ 0 ] = fresh_wire_978[ 0 ];
	assign fresh_wire_974[ 1 ] = fresh_wire_985[ 0 ];
	assign fresh_wire_974[ 2 ] = fresh_wire_986[ 0 ];
	assign fresh_wire_974[ 3 ] = fresh_wire_987[ 0 ];
	assign fresh_wire_974[ 4 ] = fresh_wire_988[ 0 ];
	assign fresh_wire_974[ 5 ] = fresh_wire_989[ 0 ];
	assign fresh_wire_974[ 6 ] = fresh_wire_990[ 0 ];
	assign fresh_wire_974[ 7 ] = fresh_wire_991[ 0 ];
	assign fresh_wire_974[ 8 ] = fresh_wire_992[ 0 ];
	assign fresh_wire_974[ 9 ] = fresh_wire_993[ 0 ];
	assign fresh_wire_974[ 10 ] = fresh_wire_979[ 0 ];
	assign fresh_wire_974[ 11 ] = fresh_wire_980[ 0 ];
	assign fresh_wire_974[ 12 ] = fresh_wire_981[ 0 ];
	assign fresh_wire_974[ 13 ] = fresh_wire_982[ 0 ];
	assign fresh_wire_974[ 14 ] = fresh_wire_983[ 0 ];
	assign fresh_wire_974[ 15 ] = fresh_wire_984[ 0 ];
	assign fresh_wire_975[ 0 ] = fresh_wire_956[ 0 ];
	assign fresh_wire_975[ 1 ] = fresh_wire_956[ 1 ];
	assign fresh_wire_975[ 2 ] = fresh_wire_956[ 2 ];
	assign fresh_wire_975[ 3 ] = fresh_wire_956[ 3 ];
	assign fresh_wire_975[ 4 ] = fresh_wire_956[ 4 ];
	assign fresh_wire_975[ 5 ] = fresh_wire_956[ 5 ];
	assign fresh_wire_975[ 6 ] = fresh_wire_956[ 6 ];
	assign fresh_wire_975[ 7 ] = fresh_wire_956[ 7 ];
	assign fresh_wire_975[ 8 ] = fresh_wire_956[ 8 ];
	assign fresh_wire_975[ 9 ] = fresh_wire_956[ 9 ];
	assign fresh_wire_975[ 10 ] = fresh_wire_956[ 10 ];
	assign fresh_wire_975[ 11 ] = fresh_wire_956[ 11 ];
	assign fresh_wire_975[ 12 ] = fresh_wire_956[ 12 ];
	assign fresh_wire_975[ 13 ] = fresh_wire_956[ 13 ];
	assign fresh_wire_975[ 14 ] = fresh_wire_956[ 14 ];
	assign fresh_wire_975[ 15 ] = fresh_wire_956[ 15 ];
	assign fresh_wire_977[ 0 ] = fresh_wire_934[ 0 ];
	assign fresh_wire_994[ 0 ] = fresh_wire_998[ 0 ];
	assign fresh_wire_994[ 1 ] = fresh_wire_999[ 0 ];
	assign fresh_wire_994[ 2 ] = fresh_wire_1000[ 0 ];
	assign fresh_wire_994[ 3 ] = fresh_wire_1001[ 0 ];
	assign fresh_wire_994[ 4 ] = fresh_wire_1002[ 0 ];
	assign fresh_wire_994[ 5 ] = fresh_wire_1003[ 0 ];
	assign fresh_wire_994[ 6 ] = fresh_wire_1004[ 0 ];
	assign fresh_wire_994[ 7 ] = fresh_wire_1005[ 0 ];
	assign fresh_wire_994[ 8 ] = fresh_wire_1006[ 0 ];
	assign fresh_wire_995[ 0 ] = fresh_wire_435[ 0 ];
	assign fresh_wire_995[ 1 ] = fresh_wire_435[ 1 ];
	assign fresh_wire_995[ 2 ] = fresh_wire_435[ 2 ];
	assign fresh_wire_995[ 3 ] = fresh_wire_435[ 3 ];
	assign fresh_wire_995[ 4 ] = fresh_wire_435[ 4 ];
	assign fresh_wire_995[ 5 ] = fresh_wire_435[ 5 ];
	assign fresh_wire_995[ 6 ] = fresh_wire_435[ 6 ];
	assign fresh_wire_995[ 7 ] = fresh_wire_435[ 7 ];
	assign fresh_wire_995[ 8 ] = fresh_wire_435[ 8 ];
	assign fresh_wire_997[ 0 ] = fresh_wire_937[ 0 ];
	assign fresh_wire_1007[ 0 ] = fresh_wire_1011[ 0 ];
	assign fresh_wire_1007[ 1 ] = fresh_wire_1012[ 0 ];
	assign fresh_wire_1007[ 2 ] = fresh_wire_1013[ 0 ];
	assign fresh_wire_1007[ 3 ] = fresh_wire_1014[ 0 ];
	assign fresh_wire_1007[ 4 ] = fresh_wire_1015[ 0 ];
	assign fresh_wire_1007[ 5 ] = fresh_wire_1016[ 0 ];
	assign fresh_wire_1007[ 6 ] = fresh_wire_1017[ 0 ];
	assign fresh_wire_1007[ 7 ] = fresh_wire_1018[ 0 ];
	assign fresh_wire_1007[ 8 ] = fresh_wire_1019[ 0 ];
	assign fresh_wire_1008[ 0 ] = fresh_wire_996[ 0 ];
	assign fresh_wire_1008[ 1 ] = fresh_wire_996[ 1 ];
	assign fresh_wire_1008[ 2 ] = fresh_wire_996[ 2 ];
	assign fresh_wire_1008[ 3 ] = fresh_wire_996[ 3 ];
	assign fresh_wire_1008[ 4 ] = fresh_wire_996[ 4 ];
	assign fresh_wire_1008[ 5 ] = fresh_wire_996[ 5 ];
	assign fresh_wire_1008[ 6 ] = fresh_wire_996[ 6 ];
	assign fresh_wire_1008[ 7 ] = fresh_wire_996[ 7 ];
	assign fresh_wire_1008[ 8 ] = fresh_wire_996[ 8 ];
	assign fresh_wire_1010[ 0 ] = fresh_wire_934[ 0 ];
	assign fresh_wire_1020[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1021[ 0 ] = fresh_wire_435[ 0 ];
	assign fresh_wire_1021[ 1 ] = fresh_wire_435[ 1 ];
	assign fresh_wire_1021[ 2 ] = fresh_wire_435[ 2 ];
	assign fresh_wire_1021[ 3 ] = fresh_wire_435[ 3 ];
	assign fresh_wire_1021[ 4 ] = fresh_wire_435[ 4 ];
	assign fresh_wire_1021[ 5 ] = fresh_wire_435[ 5 ];
	assign fresh_wire_1021[ 6 ] = fresh_wire_435[ 6 ];
	assign fresh_wire_1021[ 7 ] = fresh_wire_435[ 7 ];
	assign fresh_wire_1021[ 8 ] = fresh_wire_435[ 8 ];
	assign fresh_wire_1023[ 0 ] = fresh_wire_1009[ 0 ];
	assign fresh_wire_1023[ 1 ] = fresh_wire_1009[ 1 ];
	assign fresh_wire_1023[ 2 ] = fresh_wire_1009[ 2 ];
	assign fresh_wire_1023[ 3 ] = fresh_wire_1009[ 3 ];
	assign fresh_wire_1023[ 4 ] = fresh_wire_1009[ 4 ];
	assign fresh_wire_1023[ 5 ] = fresh_wire_1009[ 5 ];
	assign fresh_wire_1023[ 6 ] = fresh_wire_1009[ 6 ];
	assign fresh_wire_1023[ 7 ] = fresh_wire_1009[ 7 ];
	assign fresh_wire_1023[ 8 ] = fresh_wire_1009[ 8 ];
	assign fresh_wire_1024[ 0 ] = fresh_wire_976[ 0 ];
	assign fresh_wire_1024[ 1 ] = fresh_wire_976[ 1 ];
	assign fresh_wire_1024[ 2 ] = fresh_wire_976[ 2 ];
	assign fresh_wire_1024[ 3 ] = fresh_wire_976[ 3 ];
	assign fresh_wire_1024[ 4 ] = fresh_wire_976[ 4 ];
	assign fresh_wire_1024[ 5 ] = fresh_wire_976[ 5 ];
	assign fresh_wire_1024[ 6 ] = fresh_wire_976[ 6 ];
	assign fresh_wire_1024[ 7 ] = fresh_wire_976[ 7 ];
	assign fresh_wire_1024[ 8 ] = fresh_wire_976[ 8 ];
	assign fresh_wire_1024[ 9 ] = fresh_wire_976[ 9 ];
	assign fresh_wire_1024[ 10 ] = fresh_wire_976[ 10 ];
	assign fresh_wire_1024[ 11 ] = fresh_wire_976[ 11 ];
	assign fresh_wire_1024[ 12 ] = fresh_wire_976[ 12 ];
	assign fresh_wire_1024[ 13 ] = fresh_wire_976[ 13 ];
	assign fresh_wire_1024[ 14 ] = fresh_wire_976[ 14 ];
	assign fresh_wire_1024[ 15 ] = fresh_wire_976[ 15 ];
	assign fresh_wire_1025[ 0 ] = fresh_wire_952[ 0 ];
	assign fresh_wire_1026[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_1028[ 0 ] = fresh_wire_426[ 0 ];
	assign fresh_wire_1030[ 0 ] = fresh_wire_1027[ 0 ];
	assign fresh_wire_1031[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1033[ 0 ] = fresh_wire_1029[ 0 ];
	assign fresh_wire_1034[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1036[ 0 ] = fresh_wire_1041[ 0 ];
	assign fresh_wire_1036[ 1 ] = fresh_wire_1041[ 1 ];
	assign fresh_wire_1036[ 2 ] = fresh_wire_1041[ 2 ];
	assign fresh_wire_1036[ 3 ] = fresh_wire_1041[ 3 ];
	assign fresh_wire_1036[ 4 ] = fresh_wire_1041[ 4 ];
	assign fresh_wire_1036[ 5 ] = fresh_wire_1041[ 5 ];
	assign fresh_wire_1036[ 6 ] = fresh_wire_1041[ 6 ];
	assign fresh_wire_1036[ 7 ] = fresh_wire_1041[ 7 ];
	assign fresh_wire_1036[ 8 ] = fresh_wire_1041[ 8 ];
	assign fresh_wire_1036[ 9 ] = fresh_wire_1041[ 9 ];
	assign fresh_wire_1036[ 10 ] = fresh_wire_1041[ 10 ];
	assign fresh_wire_1036[ 11 ] = fresh_wire_1041[ 11 ];
	assign fresh_wire_1036[ 12 ] = fresh_wire_1041[ 12 ];
	assign fresh_wire_1036[ 13 ] = fresh_wire_1041[ 13 ];
	assign fresh_wire_1036[ 14 ] = fresh_wire_1041[ 14 ];
	assign fresh_wire_1036[ 15 ] = fresh_wire_1041[ 15 ];
	assign fresh_wire_1038[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1039[ 0 ] = fresh_wire_1037[ 0 ];
	assign fresh_wire_1039[ 1 ] = fresh_wire_1037[ 1 ];
	assign fresh_wire_1039[ 2 ] = fresh_wire_1037[ 2 ];
	assign fresh_wire_1039[ 3 ] = fresh_wire_1037[ 3 ];
	assign fresh_wire_1039[ 4 ] = fresh_wire_1037[ 4 ];
	assign fresh_wire_1039[ 5 ] = fresh_wire_1037[ 5 ];
	assign fresh_wire_1039[ 6 ] = fresh_wire_1037[ 6 ];
	assign fresh_wire_1039[ 7 ] = fresh_wire_1037[ 7 ];
	assign fresh_wire_1039[ 8 ] = fresh_wire_1037[ 8 ];
	assign fresh_wire_1039[ 9 ] = fresh_wire_1037[ 9 ];
	assign fresh_wire_1039[ 10 ] = fresh_wire_1037[ 10 ];
	assign fresh_wire_1039[ 11 ] = fresh_wire_1037[ 11 ];
	assign fresh_wire_1039[ 12 ] = fresh_wire_1037[ 12 ];
	assign fresh_wire_1039[ 13 ] = fresh_wire_1037[ 13 ];
	assign fresh_wire_1039[ 14 ] = fresh_wire_1037[ 14 ];
	assign fresh_wire_1039[ 15 ] = fresh_wire_1037[ 15 ];
	assign fresh_wire_1040[ 0 ] = fresh_wire_1120[ 0 ];
	assign fresh_wire_1040[ 1 ] = fresh_wire_1120[ 1 ];
	assign fresh_wire_1040[ 2 ] = fresh_wire_1120[ 2 ];
	assign fresh_wire_1040[ 3 ] = fresh_wire_1120[ 3 ];
	assign fresh_wire_1040[ 4 ] = fresh_wire_1120[ 4 ];
	assign fresh_wire_1040[ 5 ] = fresh_wire_1120[ 5 ];
	assign fresh_wire_1040[ 6 ] = fresh_wire_1120[ 6 ];
	assign fresh_wire_1040[ 7 ] = fresh_wire_1120[ 7 ];
	assign fresh_wire_1040[ 8 ] = fresh_wire_1120[ 8 ];
	assign fresh_wire_1040[ 9 ] = fresh_wire_1120[ 9 ];
	assign fresh_wire_1040[ 10 ] = fresh_wire_1120[ 10 ];
	assign fresh_wire_1040[ 11 ] = fresh_wire_1120[ 11 ];
	assign fresh_wire_1040[ 12 ] = fresh_wire_1120[ 12 ];
	assign fresh_wire_1040[ 13 ] = fresh_wire_1120[ 13 ];
	assign fresh_wire_1040[ 14 ] = fresh_wire_1120[ 14 ];
	assign fresh_wire_1040[ 15 ] = fresh_wire_1120[ 15 ];
	assign fresh_wire_1042[ 0 ] = fresh_wire_1032[ 0 ];
	assign fresh_wire_1043[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1043[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1043[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1043[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1043[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1043[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1043[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1043[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1043[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1043[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1043[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1043[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1043[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1043[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1043[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1043[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1044[ 0 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 1 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 2 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 3 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 4 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 5 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 6 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 7 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 8 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 9 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 10 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 11 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 12 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 13 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 14 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1044[ 15 ] = fresh_wire_1047[ 0 ];
	assign fresh_wire_1046[ 0 ] = fresh_wire_1035[ 0 ];
	assign fresh_wire_1048[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1048[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1048[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1048[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1048[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1048[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1048[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1048[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1048[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1048[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1048[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1048[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1048[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1048[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1048[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1048[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1049[ 0 ] = fresh_wire_1045[ 0 ];
	assign fresh_wire_1049[ 1 ] = fresh_wire_1045[ 1 ];
	assign fresh_wire_1049[ 2 ] = fresh_wire_1045[ 2 ];
	assign fresh_wire_1049[ 3 ] = fresh_wire_1045[ 3 ];
	assign fresh_wire_1049[ 4 ] = fresh_wire_1045[ 4 ];
	assign fresh_wire_1049[ 5 ] = fresh_wire_1045[ 5 ];
	assign fresh_wire_1049[ 6 ] = fresh_wire_1045[ 6 ];
	assign fresh_wire_1049[ 7 ] = fresh_wire_1045[ 7 ];
	assign fresh_wire_1049[ 8 ] = fresh_wire_1045[ 8 ];
	assign fresh_wire_1049[ 9 ] = fresh_wire_1045[ 9 ];
	assign fresh_wire_1049[ 10 ] = fresh_wire_1045[ 10 ];
	assign fresh_wire_1049[ 11 ] = fresh_wire_1045[ 11 ];
	assign fresh_wire_1049[ 12 ] = fresh_wire_1045[ 12 ];
	assign fresh_wire_1049[ 13 ] = fresh_wire_1045[ 13 ];
	assign fresh_wire_1049[ 14 ] = fresh_wire_1045[ 14 ];
	assign fresh_wire_1049[ 15 ] = fresh_wire_1045[ 15 ];
	assign fresh_wire_1051[ 0 ] = fresh_wire_1032[ 0 ];
	assign fresh_wire_1052[ 0 ] = fresh_wire_1056[ 0 ];
	assign fresh_wire_1052[ 1 ] = fresh_wire_1063[ 0 ];
	assign fresh_wire_1052[ 2 ] = fresh_wire_1064[ 0 ];
	assign fresh_wire_1052[ 3 ] = fresh_wire_1065[ 0 ];
	assign fresh_wire_1052[ 4 ] = fresh_wire_1066[ 0 ];
	assign fresh_wire_1052[ 5 ] = fresh_wire_1067[ 0 ];
	assign fresh_wire_1052[ 6 ] = fresh_wire_1068[ 0 ];
	assign fresh_wire_1052[ 7 ] = fresh_wire_1069[ 0 ];
	assign fresh_wire_1052[ 8 ] = fresh_wire_1070[ 0 ];
	assign fresh_wire_1052[ 9 ] = fresh_wire_1071[ 0 ];
	assign fresh_wire_1052[ 10 ] = fresh_wire_1057[ 0 ];
	assign fresh_wire_1052[ 11 ] = fresh_wire_1058[ 0 ];
	assign fresh_wire_1052[ 12 ] = fresh_wire_1059[ 0 ];
	assign fresh_wire_1052[ 13 ] = fresh_wire_1060[ 0 ];
	assign fresh_wire_1052[ 14 ] = fresh_wire_1061[ 0 ];
	assign fresh_wire_1052[ 15 ] = fresh_wire_1062[ 0 ];
	assign fresh_wire_1053[ 0 ] = fresh_wire_714[ 16 ];
	assign fresh_wire_1053[ 1 ] = fresh_wire_714[ 17 ];
	assign fresh_wire_1053[ 2 ] = fresh_wire_714[ 18 ];
	assign fresh_wire_1053[ 3 ] = fresh_wire_714[ 19 ];
	assign fresh_wire_1053[ 4 ] = fresh_wire_714[ 20 ];
	assign fresh_wire_1053[ 5 ] = fresh_wire_714[ 21 ];
	assign fresh_wire_1053[ 6 ] = fresh_wire_714[ 22 ];
	assign fresh_wire_1053[ 7 ] = fresh_wire_714[ 23 ];
	assign fresh_wire_1053[ 8 ] = fresh_wire_714[ 24 ];
	assign fresh_wire_1053[ 9 ] = fresh_wire_714[ 25 ];
	assign fresh_wire_1053[ 10 ] = fresh_wire_714[ 26 ];
	assign fresh_wire_1053[ 11 ] = fresh_wire_714[ 27 ];
	assign fresh_wire_1053[ 12 ] = fresh_wire_714[ 28 ];
	assign fresh_wire_1053[ 13 ] = fresh_wire_714[ 29 ];
	assign fresh_wire_1053[ 14 ] = fresh_wire_714[ 30 ];
	assign fresh_wire_1053[ 15 ] = fresh_wire_714[ 31 ];
	assign fresh_wire_1055[ 0 ] = fresh_wire_1035[ 0 ];
	assign fresh_wire_1072[ 0 ] = fresh_wire_1076[ 0 ];
	assign fresh_wire_1072[ 1 ] = fresh_wire_1083[ 0 ];
	assign fresh_wire_1072[ 2 ] = fresh_wire_1084[ 0 ];
	assign fresh_wire_1072[ 3 ] = fresh_wire_1085[ 0 ];
	assign fresh_wire_1072[ 4 ] = fresh_wire_1086[ 0 ];
	assign fresh_wire_1072[ 5 ] = fresh_wire_1087[ 0 ];
	assign fresh_wire_1072[ 6 ] = fresh_wire_1088[ 0 ];
	assign fresh_wire_1072[ 7 ] = fresh_wire_1089[ 0 ];
	assign fresh_wire_1072[ 8 ] = fresh_wire_1090[ 0 ];
	assign fresh_wire_1072[ 9 ] = fresh_wire_1091[ 0 ];
	assign fresh_wire_1072[ 10 ] = fresh_wire_1077[ 0 ];
	assign fresh_wire_1072[ 11 ] = fresh_wire_1078[ 0 ];
	assign fresh_wire_1072[ 12 ] = fresh_wire_1079[ 0 ];
	assign fresh_wire_1072[ 13 ] = fresh_wire_1080[ 0 ];
	assign fresh_wire_1072[ 14 ] = fresh_wire_1081[ 0 ];
	assign fresh_wire_1072[ 15 ] = fresh_wire_1082[ 0 ];
	assign fresh_wire_1073[ 0 ] = fresh_wire_1054[ 0 ];
	assign fresh_wire_1073[ 1 ] = fresh_wire_1054[ 1 ];
	assign fresh_wire_1073[ 2 ] = fresh_wire_1054[ 2 ];
	assign fresh_wire_1073[ 3 ] = fresh_wire_1054[ 3 ];
	assign fresh_wire_1073[ 4 ] = fresh_wire_1054[ 4 ];
	assign fresh_wire_1073[ 5 ] = fresh_wire_1054[ 5 ];
	assign fresh_wire_1073[ 6 ] = fresh_wire_1054[ 6 ];
	assign fresh_wire_1073[ 7 ] = fresh_wire_1054[ 7 ];
	assign fresh_wire_1073[ 8 ] = fresh_wire_1054[ 8 ];
	assign fresh_wire_1073[ 9 ] = fresh_wire_1054[ 9 ];
	assign fresh_wire_1073[ 10 ] = fresh_wire_1054[ 10 ];
	assign fresh_wire_1073[ 11 ] = fresh_wire_1054[ 11 ];
	assign fresh_wire_1073[ 12 ] = fresh_wire_1054[ 12 ];
	assign fresh_wire_1073[ 13 ] = fresh_wire_1054[ 13 ];
	assign fresh_wire_1073[ 14 ] = fresh_wire_1054[ 14 ];
	assign fresh_wire_1073[ 15 ] = fresh_wire_1054[ 15 ];
	assign fresh_wire_1075[ 0 ] = fresh_wire_1032[ 0 ];
	assign fresh_wire_1092[ 0 ] = fresh_wire_1096[ 0 ];
	assign fresh_wire_1092[ 1 ] = fresh_wire_1097[ 0 ];
	assign fresh_wire_1092[ 2 ] = fresh_wire_1098[ 0 ];
	assign fresh_wire_1092[ 3 ] = fresh_wire_1099[ 0 ];
	assign fresh_wire_1092[ 4 ] = fresh_wire_1100[ 0 ];
	assign fresh_wire_1092[ 5 ] = fresh_wire_1101[ 0 ];
	assign fresh_wire_1092[ 6 ] = fresh_wire_1102[ 0 ];
	assign fresh_wire_1092[ 7 ] = fresh_wire_1103[ 0 ];
	assign fresh_wire_1092[ 8 ] = fresh_wire_1104[ 0 ];
	assign fresh_wire_1093[ 0 ] = fresh_wire_435[ 0 ];
	assign fresh_wire_1093[ 1 ] = fresh_wire_435[ 1 ];
	assign fresh_wire_1093[ 2 ] = fresh_wire_435[ 2 ];
	assign fresh_wire_1093[ 3 ] = fresh_wire_435[ 3 ];
	assign fresh_wire_1093[ 4 ] = fresh_wire_435[ 4 ];
	assign fresh_wire_1093[ 5 ] = fresh_wire_435[ 5 ];
	assign fresh_wire_1093[ 6 ] = fresh_wire_435[ 6 ];
	assign fresh_wire_1093[ 7 ] = fresh_wire_435[ 7 ];
	assign fresh_wire_1093[ 8 ] = fresh_wire_435[ 8 ];
	assign fresh_wire_1095[ 0 ] = fresh_wire_1035[ 0 ];
	assign fresh_wire_1105[ 0 ] = fresh_wire_1109[ 0 ];
	assign fresh_wire_1105[ 1 ] = fresh_wire_1110[ 0 ];
	assign fresh_wire_1105[ 2 ] = fresh_wire_1111[ 0 ];
	assign fresh_wire_1105[ 3 ] = fresh_wire_1112[ 0 ];
	assign fresh_wire_1105[ 4 ] = fresh_wire_1113[ 0 ];
	assign fresh_wire_1105[ 5 ] = fresh_wire_1114[ 0 ];
	assign fresh_wire_1105[ 6 ] = fresh_wire_1115[ 0 ];
	assign fresh_wire_1105[ 7 ] = fresh_wire_1116[ 0 ];
	assign fresh_wire_1105[ 8 ] = fresh_wire_1117[ 0 ];
	assign fresh_wire_1106[ 0 ] = fresh_wire_1094[ 0 ];
	assign fresh_wire_1106[ 1 ] = fresh_wire_1094[ 1 ];
	assign fresh_wire_1106[ 2 ] = fresh_wire_1094[ 2 ];
	assign fresh_wire_1106[ 3 ] = fresh_wire_1094[ 3 ];
	assign fresh_wire_1106[ 4 ] = fresh_wire_1094[ 4 ];
	assign fresh_wire_1106[ 5 ] = fresh_wire_1094[ 5 ];
	assign fresh_wire_1106[ 6 ] = fresh_wire_1094[ 6 ];
	assign fresh_wire_1106[ 7 ] = fresh_wire_1094[ 7 ];
	assign fresh_wire_1106[ 8 ] = fresh_wire_1094[ 8 ];
	assign fresh_wire_1108[ 0 ] = fresh_wire_1032[ 0 ];
	assign fresh_wire_1118[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1119[ 0 ] = fresh_wire_435[ 0 ];
	assign fresh_wire_1119[ 1 ] = fresh_wire_435[ 1 ];
	assign fresh_wire_1119[ 2 ] = fresh_wire_435[ 2 ];
	assign fresh_wire_1119[ 3 ] = fresh_wire_435[ 3 ];
	assign fresh_wire_1119[ 4 ] = fresh_wire_435[ 4 ];
	assign fresh_wire_1119[ 5 ] = fresh_wire_435[ 5 ];
	assign fresh_wire_1119[ 6 ] = fresh_wire_435[ 6 ];
	assign fresh_wire_1119[ 7 ] = fresh_wire_435[ 7 ];
	assign fresh_wire_1119[ 8 ] = fresh_wire_435[ 8 ];
	assign fresh_wire_1121[ 0 ] = fresh_wire_1107[ 0 ];
	assign fresh_wire_1121[ 1 ] = fresh_wire_1107[ 1 ];
	assign fresh_wire_1121[ 2 ] = fresh_wire_1107[ 2 ];
	assign fresh_wire_1121[ 3 ] = fresh_wire_1107[ 3 ];
	assign fresh_wire_1121[ 4 ] = fresh_wire_1107[ 4 ];
	assign fresh_wire_1121[ 5 ] = fresh_wire_1107[ 5 ];
	assign fresh_wire_1121[ 6 ] = fresh_wire_1107[ 6 ];
	assign fresh_wire_1121[ 7 ] = fresh_wire_1107[ 7 ];
	assign fresh_wire_1121[ 8 ] = fresh_wire_1107[ 8 ];
	assign fresh_wire_1122[ 0 ] = fresh_wire_1074[ 0 ];
	assign fresh_wire_1122[ 1 ] = fresh_wire_1074[ 1 ];
	assign fresh_wire_1122[ 2 ] = fresh_wire_1074[ 2 ];
	assign fresh_wire_1122[ 3 ] = fresh_wire_1074[ 3 ];
	assign fresh_wire_1122[ 4 ] = fresh_wire_1074[ 4 ];
	assign fresh_wire_1122[ 5 ] = fresh_wire_1074[ 5 ];
	assign fresh_wire_1122[ 6 ] = fresh_wire_1074[ 6 ];
	assign fresh_wire_1122[ 7 ] = fresh_wire_1074[ 7 ];
	assign fresh_wire_1122[ 8 ] = fresh_wire_1074[ 8 ];
	assign fresh_wire_1122[ 9 ] = fresh_wire_1074[ 9 ];
	assign fresh_wire_1122[ 10 ] = fresh_wire_1074[ 10 ];
	assign fresh_wire_1122[ 11 ] = fresh_wire_1074[ 11 ];
	assign fresh_wire_1122[ 12 ] = fresh_wire_1074[ 12 ];
	assign fresh_wire_1122[ 13 ] = fresh_wire_1074[ 13 ];
	assign fresh_wire_1122[ 14 ] = fresh_wire_1074[ 14 ];
	assign fresh_wire_1122[ 15 ] = fresh_wire_1074[ 15 ];
	assign fresh_wire_1123[ 0 ] = fresh_wire_1050[ 0 ];
	assign fresh_wire_1124[ 0 ] = fresh_wire_609[ 0 ];
	assign fresh_wire_1124[ 1 ] = fresh_wire_609[ 1 ];
	assign fresh_wire_1124[ 2 ] = fresh_wire_609[ 2 ];
	assign fresh_wire_1124[ 3 ] = fresh_wire_609[ 3 ];
	assign fresh_wire_1124[ 4 ] = fresh_wire_609[ 4 ];
	assign fresh_wire_1124[ 5 ] = fresh_wire_609[ 5 ];
	assign fresh_wire_1124[ 6 ] = fresh_wire_609[ 6 ];
	assign fresh_wire_1124[ 7 ] = fresh_wire_609[ 7 ];
	assign fresh_wire_1124[ 8 ] = fresh_wire_609[ 8 ];
	assign fresh_wire_1124[ 9 ] = fresh_wire_609[ 9 ];
	assign fresh_wire_1124[ 10 ] = fresh_wire_609[ 10 ];
	assign fresh_wire_1124[ 11 ] = fresh_wire_609[ 11 ];
	assign fresh_wire_1124[ 12 ] = fresh_wire_609[ 12 ];
	assign fresh_wire_1124[ 13 ] = fresh_wire_609[ 13 ];
	assign fresh_wire_1124[ 14 ] = fresh_wire_609[ 14 ];
	assign fresh_wire_1124[ 15 ] = fresh_wire_609[ 15 ];
	assign fresh_wire_1126[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1127[ 0 ] = fresh_wire_2177[ 0 ];
	assign fresh_wire_1128[ 0 ] = fresh_wire_1135[ 0 ];
	assign fresh_wire_1130[ 0 ] = fresh_wire_2177[ 0 ];
	assign fresh_wire_1131[ 0 ] = fresh_wire_1135[ 0 ];
	assign fresh_wire_1133[ 0 ] = fresh_wire_1398[ 0 ];
	assign fresh_wire_1134[ 0 ] = fresh_wire_1173[ 0 ];
	assign fresh_wire_1136[ 0 ] = fresh_wire_1378[ 0 ];
	assign fresh_wire_1136[ 1 ] = fresh_wire_1378[ 1 ];
	assign fresh_wire_1136[ 2 ] = fresh_wire_1378[ 2 ];
	assign fresh_wire_1136[ 3 ] = fresh_wire_1378[ 3 ];
	assign fresh_wire_1136[ 4 ] = fresh_wire_1378[ 4 ];
	assign fresh_wire_1136[ 5 ] = fresh_wire_1378[ 5 ];
	assign fresh_wire_1136[ 6 ] = fresh_wire_1378[ 6 ];
	assign fresh_wire_1136[ 7 ] = fresh_wire_1378[ 7 ];
	assign fresh_wire_1136[ 8 ] = fresh_wire_1378[ 8 ];
	assign fresh_wire_1136[ 9 ] = fresh_wire_1378[ 9 ];
	assign fresh_wire_1136[ 10 ] = fresh_wire_1378[ 10 ];
	assign fresh_wire_1136[ 11 ] = fresh_wire_1378[ 11 ];
	assign fresh_wire_1136[ 12 ] = fresh_wire_1378[ 12 ];
	assign fresh_wire_1136[ 13 ] = fresh_wire_1378[ 13 ];
	assign fresh_wire_1136[ 14 ] = fresh_wire_1378[ 14 ];
	assign fresh_wire_1136[ 15 ] = fresh_wire_1378[ 15 ];
	assign fresh_wire_1137[ 0 ] = fresh_wire_2260[ 0 ];
	assign fresh_wire_1137[ 1 ] = fresh_wire_2260[ 1 ];
	assign fresh_wire_1137[ 2 ] = fresh_wire_2260[ 2 ];
	assign fresh_wire_1137[ 3 ] = fresh_wire_2260[ 3 ];
	assign fresh_wire_1137[ 4 ] = fresh_wire_2260[ 4 ];
	assign fresh_wire_1137[ 5 ] = fresh_wire_2260[ 5 ];
	assign fresh_wire_1137[ 6 ] = fresh_wire_2260[ 6 ];
	assign fresh_wire_1137[ 7 ] = fresh_wire_2260[ 7 ];
	assign fresh_wire_1137[ 8 ] = fresh_wire_2260[ 8 ];
	assign fresh_wire_1137[ 9 ] = fresh_wire_2260[ 9 ];
	assign fresh_wire_1137[ 10 ] = fresh_wire_2260[ 10 ];
	assign fresh_wire_1137[ 11 ] = fresh_wire_2260[ 11 ];
	assign fresh_wire_1137[ 12 ] = fresh_wire_2260[ 12 ];
	assign fresh_wire_1137[ 13 ] = fresh_wire_2260[ 13 ];
	assign fresh_wire_1137[ 14 ] = fresh_wire_2260[ 14 ];
	assign fresh_wire_1137[ 15 ] = fresh_wire_2260[ 15 ];
	assign fresh_wire_1139[ 0 ] = fresh_wire_1638[ 0 ];
	assign fresh_wire_1139[ 1 ] = fresh_wire_1638[ 1 ];
	assign fresh_wire_1141[ 0 ] = fresh_wire_1390[ 0 ];
	assign fresh_wire_1141[ 1 ] = fresh_wire_1390[ 1 ];
	assign fresh_wire_1141[ 2 ] = fresh_wire_1390[ 2 ];
	assign fresh_wire_1141[ 3 ] = fresh_wire_1390[ 3 ];
	assign fresh_wire_1141[ 4 ] = fresh_wire_1390[ 4 ];
	assign fresh_wire_1141[ 5 ] = fresh_wire_1390[ 5 ];
	assign fresh_wire_1141[ 6 ] = fresh_wire_1390[ 6 ];
	assign fresh_wire_1141[ 7 ] = fresh_wire_1390[ 7 ];
	assign fresh_wire_1141[ 8 ] = fresh_wire_1390[ 8 ];
	assign fresh_wire_1141[ 9 ] = fresh_wire_1390[ 9 ];
	assign fresh_wire_1141[ 10 ] = fresh_wire_1390[ 10 ];
	assign fresh_wire_1141[ 11 ] = fresh_wire_1390[ 11 ];
	assign fresh_wire_1141[ 12 ] = fresh_wire_1390[ 12 ];
	assign fresh_wire_1141[ 13 ] = fresh_wire_1390[ 13 ];
	assign fresh_wire_1141[ 14 ] = fresh_wire_1390[ 14 ];
	assign fresh_wire_1141[ 15 ] = fresh_wire_1390[ 15 ];
	assign fresh_wire_1142[ 0 ] = fresh_wire_1140[ 0 ];
	assign fresh_wire_1142[ 1 ] = fresh_wire_1140[ 1 ];
	assign fresh_wire_1142[ 2 ] = fresh_wire_1140[ 2 ];
	assign fresh_wire_1142[ 3 ] = fresh_wire_1140[ 3 ];
	assign fresh_wire_1142[ 4 ] = fresh_wire_1140[ 4 ];
	assign fresh_wire_1142[ 5 ] = fresh_wire_1140[ 5 ];
	assign fresh_wire_1142[ 6 ] = fresh_wire_1140[ 6 ];
	assign fresh_wire_1142[ 7 ] = fresh_wire_1140[ 7 ];
	assign fresh_wire_1142[ 8 ] = fresh_wire_1140[ 8 ];
	assign fresh_wire_1142[ 9 ] = fresh_wire_1140[ 9 ];
	assign fresh_wire_1142[ 10 ] = fresh_wire_1140[ 10 ];
	assign fresh_wire_1142[ 11 ] = fresh_wire_1140[ 11 ];
	assign fresh_wire_1142[ 12 ] = fresh_wire_1140[ 12 ];
	assign fresh_wire_1142[ 13 ] = fresh_wire_1140[ 13 ];
	assign fresh_wire_1142[ 14 ] = fresh_wire_1140[ 14 ];
	assign fresh_wire_1142[ 15 ] = fresh_wire_1140[ 15 ];
	assign fresh_wire_1144[ 0 ] = fresh_wire_1386[ 0 ];
	assign fresh_wire_1144[ 1 ] = fresh_wire_1386[ 1 ];
	assign fresh_wire_1144[ 2 ] = fresh_wire_1386[ 2 ];
	assign fresh_wire_1144[ 3 ] = fresh_wire_1386[ 3 ];
	assign fresh_wire_1144[ 4 ] = fresh_wire_1386[ 4 ];
	assign fresh_wire_1144[ 5 ] = fresh_wire_1386[ 5 ];
	assign fresh_wire_1144[ 6 ] = fresh_wire_1386[ 6 ];
	assign fresh_wire_1144[ 7 ] = fresh_wire_1386[ 7 ];
	assign fresh_wire_1144[ 8 ] = fresh_wire_1386[ 8 ];
	assign fresh_wire_1144[ 9 ] = fresh_wire_1386[ 9 ];
	assign fresh_wire_1144[ 10 ] = fresh_wire_1386[ 10 ];
	assign fresh_wire_1144[ 11 ] = fresh_wire_1386[ 11 ];
	assign fresh_wire_1144[ 12 ] = fresh_wire_1386[ 12 ];
	assign fresh_wire_1144[ 13 ] = fresh_wire_1386[ 13 ];
	assign fresh_wire_1144[ 14 ] = fresh_wire_1386[ 14 ];
	assign fresh_wire_1144[ 15 ] = fresh_wire_1386[ 15 ];
	assign fresh_wire_1146[ 0 ] = fresh_wire_1145[ 0 ];
	assign fresh_wire_1146[ 1 ] = fresh_wire_1145[ 1 ];
	assign fresh_wire_1146[ 2 ] = fresh_wire_1145[ 2 ];
	assign fresh_wire_1146[ 3 ] = fresh_wire_1145[ 3 ];
	assign fresh_wire_1146[ 4 ] = fresh_wire_1145[ 4 ];
	assign fresh_wire_1146[ 5 ] = fresh_wire_1145[ 5 ];
	assign fresh_wire_1146[ 6 ] = fresh_wire_1145[ 6 ];
	assign fresh_wire_1146[ 7 ] = fresh_wire_1145[ 7 ];
	assign fresh_wire_1146[ 8 ] = fresh_wire_1145[ 8 ];
	assign fresh_wire_1146[ 9 ] = fresh_wire_1145[ 9 ];
	assign fresh_wire_1146[ 10 ] = fresh_wire_1145[ 10 ];
	assign fresh_wire_1146[ 11 ] = fresh_wire_1145[ 11 ];
	assign fresh_wire_1146[ 12 ] = fresh_wire_1145[ 12 ];
	assign fresh_wire_1146[ 13 ] = fresh_wire_1145[ 13 ];
	assign fresh_wire_1146[ 14 ] = fresh_wire_1145[ 14 ];
	assign fresh_wire_1146[ 15 ] = fresh_wire_1145[ 15 ];
	assign fresh_wire_1146[ 16 ] = fresh_wire_1145[ 16 ];
	assign fresh_wire_1146[ 17 ] = fresh_wire_1145[ 17 ];
	assign fresh_wire_1146[ 18 ] = fresh_wire_1145[ 18 ];
	assign fresh_wire_1146[ 19 ] = fresh_wire_1145[ 19 ];
	assign fresh_wire_1146[ 20 ] = fresh_wire_1145[ 20 ];
	assign fresh_wire_1146[ 21 ] = fresh_wire_1145[ 21 ];
	assign fresh_wire_1146[ 22 ] = fresh_wire_1145[ 22 ];
	assign fresh_wire_1146[ 23 ] = fresh_wire_1145[ 23 ];
	assign fresh_wire_1146[ 24 ] = fresh_wire_1145[ 24 ];
	assign fresh_wire_1146[ 25 ] = fresh_wire_1145[ 25 ];
	assign fresh_wire_1146[ 26 ] = fresh_wire_1145[ 26 ];
	assign fresh_wire_1146[ 27 ] = fresh_wire_1145[ 27 ];
	assign fresh_wire_1146[ 28 ] = fresh_wire_1145[ 28 ];
	assign fresh_wire_1146[ 29 ] = fresh_wire_1145[ 29 ];
	assign fresh_wire_1146[ 30 ] = fresh_wire_1145[ 30 ];
	assign fresh_wire_1146[ 31 ] = fresh_wire_1145[ 31 ];
	assign fresh_wire_1147[ 0 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1147[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 16 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 17 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 18 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 19 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 20 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 21 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 22 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 23 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 24 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 25 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 26 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 27 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 28 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 29 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 30 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1147[ 31 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1149[ 0 ] = fresh_wire_1390[ 0 ];
	assign fresh_wire_1149[ 1 ] = fresh_wire_1390[ 1 ];
	assign fresh_wire_1149[ 2 ] = fresh_wire_1390[ 2 ];
	assign fresh_wire_1149[ 3 ] = fresh_wire_1390[ 3 ];
	assign fresh_wire_1149[ 4 ] = fresh_wire_1390[ 4 ];
	assign fresh_wire_1149[ 5 ] = fresh_wire_1390[ 5 ];
	assign fresh_wire_1149[ 6 ] = fresh_wire_1390[ 6 ];
	assign fresh_wire_1149[ 7 ] = fresh_wire_1390[ 7 ];
	assign fresh_wire_1149[ 8 ] = fresh_wire_1390[ 8 ];
	assign fresh_wire_1149[ 9 ] = fresh_wire_1390[ 9 ];
	assign fresh_wire_1149[ 10 ] = fresh_wire_1390[ 10 ];
	assign fresh_wire_1149[ 11 ] = fresh_wire_1390[ 11 ];
	assign fresh_wire_1149[ 12 ] = fresh_wire_1390[ 12 ];
	assign fresh_wire_1149[ 13 ] = fresh_wire_1390[ 13 ];
	assign fresh_wire_1149[ 14 ] = fresh_wire_1390[ 14 ];
	assign fresh_wire_1149[ 15 ] = fresh_wire_1390[ 15 ];
	assign fresh_wire_1151[ 0 ] = fresh_wire_1150[ 0 ];
	assign fresh_wire_1151[ 1 ] = fresh_wire_1150[ 1 ];
	assign fresh_wire_1151[ 2 ] = fresh_wire_1150[ 2 ];
	assign fresh_wire_1151[ 3 ] = fresh_wire_1150[ 3 ];
	assign fresh_wire_1151[ 4 ] = fresh_wire_1150[ 4 ];
	assign fresh_wire_1151[ 5 ] = fresh_wire_1150[ 5 ];
	assign fresh_wire_1151[ 6 ] = fresh_wire_1150[ 6 ];
	assign fresh_wire_1151[ 7 ] = fresh_wire_1150[ 7 ];
	assign fresh_wire_1151[ 8 ] = fresh_wire_1150[ 8 ];
	assign fresh_wire_1151[ 9 ] = fresh_wire_1150[ 9 ];
	assign fresh_wire_1151[ 10 ] = fresh_wire_1150[ 10 ];
	assign fresh_wire_1151[ 11 ] = fresh_wire_1150[ 11 ];
	assign fresh_wire_1151[ 12 ] = fresh_wire_1150[ 12 ];
	assign fresh_wire_1151[ 13 ] = fresh_wire_1150[ 13 ];
	assign fresh_wire_1151[ 14 ] = fresh_wire_1150[ 14 ];
	assign fresh_wire_1151[ 15 ] = fresh_wire_1150[ 15 ];
	assign fresh_wire_1151[ 16 ] = fresh_wire_1150[ 16 ];
	assign fresh_wire_1151[ 17 ] = fresh_wire_1150[ 17 ];
	assign fresh_wire_1151[ 18 ] = fresh_wire_1150[ 18 ];
	assign fresh_wire_1151[ 19 ] = fresh_wire_1150[ 19 ];
	assign fresh_wire_1151[ 20 ] = fresh_wire_1150[ 20 ];
	assign fresh_wire_1151[ 21 ] = fresh_wire_1150[ 21 ];
	assign fresh_wire_1151[ 22 ] = fresh_wire_1150[ 22 ];
	assign fresh_wire_1151[ 23 ] = fresh_wire_1150[ 23 ];
	assign fresh_wire_1151[ 24 ] = fresh_wire_1150[ 24 ];
	assign fresh_wire_1151[ 25 ] = fresh_wire_1150[ 25 ];
	assign fresh_wire_1151[ 26 ] = fresh_wire_1150[ 26 ];
	assign fresh_wire_1151[ 27 ] = fresh_wire_1150[ 27 ];
	assign fresh_wire_1151[ 28 ] = fresh_wire_1150[ 28 ];
	assign fresh_wire_1151[ 29 ] = fresh_wire_1150[ 29 ];
	assign fresh_wire_1151[ 30 ] = fresh_wire_1150[ 30 ];
	assign fresh_wire_1151[ 31 ] = fresh_wire_1150[ 31 ];
	assign fresh_wire_1152[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 1 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1152[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 16 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 17 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 18 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 19 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 20 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 21 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 22 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 23 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 24 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 25 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 26 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 27 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 28 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 29 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 30 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1152[ 31 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1154[ 0 ] = fresh_wire_1382[ 0 ];
	assign fresh_wire_1154[ 1 ] = fresh_wire_1382[ 1 ];
	assign fresh_wire_1154[ 2 ] = fresh_wire_1382[ 2 ];
	assign fresh_wire_1154[ 3 ] = fresh_wire_1382[ 3 ];
	assign fresh_wire_1154[ 4 ] = fresh_wire_1382[ 4 ];
	assign fresh_wire_1154[ 5 ] = fresh_wire_1382[ 5 ];
	assign fresh_wire_1154[ 6 ] = fresh_wire_1382[ 6 ];
	assign fresh_wire_1154[ 7 ] = fresh_wire_1382[ 7 ];
	assign fresh_wire_1154[ 8 ] = fresh_wire_1382[ 8 ];
	assign fresh_wire_1154[ 9 ] = fresh_wire_1382[ 9 ];
	assign fresh_wire_1154[ 10 ] = fresh_wire_1382[ 10 ];
	assign fresh_wire_1154[ 11 ] = fresh_wire_1382[ 11 ];
	assign fresh_wire_1154[ 12 ] = fresh_wire_1382[ 12 ];
	assign fresh_wire_1154[ 13 ] = fresh_wire_1382[ 13 ];
	assign fresh_wire_1154[ 14 ] = fresh_wire_1382[ 14 ];
	assign fresh_wire_1154[ 15 ] = fresh_wire_1382[ 15 ];
	assign fresh_wire_1156[ 0 ] = fresh_wire_1155[ 0 ];
	assign fresh_wire_1156[ 1 ] = fresh_wire_1155[ 1 ];
	assign fresh_wire_1156[ 2 ] = fresh_wire_1155[ 2 ];
	assign fresh_wire_1156[ 3 ] = fresh_wire_1155[ 3 ];
	assign fresh_wire_1156[ 4 ] = fresh_wire_1155[ 4 ];
	assign fresh_wire_1156[ 5 ] = fresh_wire_1155[ 5 ];
	assign fresh_wire_1156[ 6 ] = fresh_wire_1155[ 6 ];
	assign fresh_wire_1156[ 7 ] = fresh_wire_1155[ 7 ];
	assign fresh_wire_1156[ 8 ] = fresh_wire_1155[ 8 ];
	assign fresh_wire_1156[ 9 ] = fresh_wire_1155[ 9 ];
	assign fresh_wire_1156[ 10 ] = fresh_wire_1155[ 10 ];
	assign fresh_wire_1156[ 11 ] = fresh_wire_1155[ 11 ];
	assign fresh_wire_1156[ 12 ] = fresh_wire_1155[ 12 ];
	assign fresh_wire_1156[ 13 ] = fresh_wire_1155[ 13 ];
	assign fresh_wire_1156[ 14 ] = fresh_wire_1155[ 14 ];
	assign fresh_wire_1156[ 15 ] = fresh_wire_1155[ 15 ];
	assign fresh_wire_1156[ 16 ] = fresh_wire_1155[ 16 ];
	assign fresh_wire_1156[ 17 ] = fresh_wire_1155[ 17 ];
	assign fresh_wire_1156[ 18 ] = fresh_wire_1155[ 18 ];
	assign fresh_wire_1156[ 19 ] = fresh_wire_1155[ 19 ];
	assign fresh_wire_1156[ 20 ] = fresh_wire_1155[ 20 ];
	assign fresh_wire_1156[ 21 ] = fresh_wire_1155[ 21 ];
	assign fresh_wire_1156[ 22 ] = fresh_wire_1155[ 22 ];
	assign fresh_wire_1156[ 23 ] = fresh_wire_1155[ 23 ];
	assign fresh_wire_1156[ 24 ] = fresh_wire_1155[ 24 ];
	assign fresh_wire_1156[ 25 ] = fresh_wire_1155[ 25 ];
	assign fresh_wire_1156[ 26 ] = fresh_wire_1155[ 26 ];
	assign fresh_wire_1156[ 27 ] = fresh_wire_1155[ 27 ];
	assign fresh_wire_1156[ 28 ] = fresh_wire_1155[ 28 ];
	assign fresh_wire_1156[ 29 ] = fresh_wire_1155[ 29 ];
	assign fresh_wire_1156[ 30 ] = fresh_wire_1155[ 30 ];
	assign fresh_wire_1156[ 31 ] = fresh_wire_1155[ 31 ];
	assign fresh_wire_1157[ 0 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1157[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 16 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 17 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 18 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 19 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 20 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 21 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 22 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 23 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 24 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 25 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 26 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 27 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 28 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 29 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 30 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1157[ 31 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1159[ 0 ] = fresh_wire_1378[ 0 ];
	assign fresh_wire_1159[ 1 ] = fresh_wire_1378[ 1 ];
	assign fresh_wire_1159[ 2 ] = fresh_wire_1378[ 2 ];
	assign fresh_wire_1159[ 3 ] = fresh_wire_1378[ 3 ];
	assign fresh_wire_1159[ 4 ] = fresh_wire_1378[ 4 ];
	assign fresh_wire_1159[ 5 ] = fresh_wire_1378[ 5 ];
	assign fresh_wire_1159[ 6 ] = fresh_wire_1378[ 6 ];
	assign fresh_wire_1159[ 7 ] = fresh_wire_1378[ 7 ];
	assign fresh_wire_1159[ 8 ] = fresh_wire_1378[ 8 ];
	assign fresh_wire_1159[ 9 ] = fresh_wire_1378[ 9 ];
	assign fresh_wire_1159[ 10 ] = fresh_wire_1378[ 10 ];
	assign fresh_wire_1159[ 11 ] = fresh_wire_1378[ 11 ];
	assign fresh_wire_1159[ 12 ] = fresh_wire_1378[ 12 ];
	assign fresh_wire_1159[ 13 ] = fresh_wire_1378[ 13 ];
	assign fresh_wire_1159[ 14 ] = fresh_wire_1378[ 14 ];
	assign fresh_wire_1159[ 15 ] = fresh_wire_1378[ 15 ];
	assign fresh_wire_1160[ 0 ] = fresh_wire_2261[ 0 ];
	assign fresh_wire_1160[ 1 ] = fresh_wire_2261[ 1 ];
	assign fresh_wire_1160[ 2 ] = fresh_wire_2261[ 2 ];
	assign fresh_wire_1160[ 3 ] = fresh_wire_2261[ 3 ];
	assign fresh_wire_1160[ 4 ] = fresh_wire_2261[ 4 ];
	assign fresh_wire_1160[ 5 ] = fresh_wire_2261[ 5 ];
	assign fresh_wire_1160[ 6 ] = fresh_wire_2261[ 6 ];
	assign fresh_wire_1160[ 7 ] = fresh_wire_2261[ 7 ];
	assign fresh_wire_1160[ 8 ] = fresh_wire_2261[ 8 ];
	assign fresh_wire_1160[ 9 ] = fresh_wire_2261[ 9 ];
	assign fresh_wire_1160[ 10 ] = fresh_wire_2261[ 10 ];
	assign fresh_wire_1160[ 11 ] = fresh_wire_2261[ 11 ];
	assign fresh_wire_1160[ 12 ] = fresh_wire_2261[ 12 ];
	assign fresh_wire_1160[ 13 ] = fresh_wire_2261[ 13 ];
	assign fresh_wire_1160[ 14 ] = fresh_wire_2261[ 14 ];
	assign fresh_wire_1160[ 15 ] = fresh_wire_2261[ 15 ];
	assign fresh_wire_1162[ 0 ] = fresh_wire_1378[ 0 ];
	assign fresh_wire_1162[ 1 ] = fresh_wire_1378[ 1 ];
	assign fresh_wire_1162[ 2 ] = fresh_wire_1378[ 2 ];
	assign fresh_wire_1162[ 3 ] = fresh_wire_1378[ 3 ];
	assign fresh_wire_1162[ 4 ] = fresh_wire_1378[ 4 ];
	assign fresh_wire_1162[ 5 ] = fresh_wire_1378[ 5 ];
	assign fresh_wire_1162[ 6 ] = fresh_wire_1378[ 6 ];
	assign fresh_wire_1162[ 7 ] = fresh_wire_1378[ 7 ];
	assign fresh_wire_1162[ 8 ] = fresh_wire_1378[ 8 ];
	assign fresh_wire_1162[ 9 ] = fresh_wire_1378[ 9 ];
	assign fresh_wire_1162[ 10 ] = fresh_wire_1378[ 10 ];
	assign fresh_wire_1162[ 11 ] = fresh_wire_1378[ 11 ];
	assign fresh_wire_1162[ 12 ] = fresh_wire_1378[ 12 ];
	assign fresh_wire_1162[ 13 ] = fresh_wire_1378[ 13 ];
	assign fresh_wire_1162[ 14 ] = fresh_wire_1378[ 14 ];
	assign fresh_wire_1162[ 15 ] = fresh_wire_1378[ 15 ];
	assign fresh_wire_1163[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1163[ 1 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1163[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1163[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1163[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1163[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1163[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1163[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1163[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1163[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1163[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1163[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1163[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1163[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1163[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1163[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1165[ 0 ] = fresh_wire_1378[ 0 ];
	assign fresh_wire_1165[ 1 ] = fresh_wire_1378[ 1 ];
	assign fresh_wire_1165[ 2 ] = fresh_wire_1378[ 2 ];
	assign fresh_wire_1165[ 3 ] = fresh_wire_1378[ 3 ];
	assign fresh_wire_1165[ 4 ] = fresh_wire_1378[ 4 ];
	assign fresh_wire_1165[ 5 ] = fresh_wire_1378[ 5 ];
	assign fresh_wire_1165[ 6 ] = fresh_wire_1378[ 6 ];
	assign fresh_wire_1165[ 7 ] = fresh_wire_1378[ 7 ];
	assign fresh_wire_1165[ 8 ] = fresh_wire_1378[ 8 ];
	assign fresh_wire_1165[ 9 ] = fresh_wire_1378[ 9 ];
	assign fresh_wire_1165[ 10 ] = fresh_wire_1378[ 10 ];
	assign fresh_wire_1165[ 11 ] = fresh_wire_1378[ 11 ];
	assign fresh_wire_1165[ 12 ] = fresh_wire_1378[ 12 ];
	assign fresh_wire_1165[ 13 ] = fresh_wire_1378[ 13 ];
	assign fresh_wire_1165[ 14 ] = fresh_wire_1378[ 14 ];
	assign fresh_wire_1165[ 15 ] = fresh_wire_1378[ 15 ];
	assign fresh_wire_1166[ 0 ] = fresh_wire_2262[ 0 ];
	assign fresh_wire_1166[ 1 ] = fresh_wire_2262[ 1 ];
	assign fresh_wire_1166[ 2 ] = fresh_wire_2262[ 2 ];
	assign fresh_wire_1166[ 3 ] = fresh_wire_2262[ 3 ];
	assign fresh_wire_1166[ 4 ] = fresh_wire_2262[ 4 ];
	assign fresh_wire_1166[ 5 ] = fresh_wire_2262[ 5 ];
	assign fresh_wire_1166[ 6 ] = fresh_wire_2262[ 6 ];
	assign fresh_wire_1166[ 7 ] = fresh_wire_2262[ 7 ];
	assign fresh_wire_1166[ 8 ] = fresh_wire_2262[ 8 ];
	assign fresh_wire_1166[ 9 ] = fresh_wire_2262[ 9 ];
	assign fresh_wire_1166[ 10 ] = fresh_wire_2262[ 10 ];
	assign fresh_wire_1166[ 11 ] = fresh_wire_2262[ 11 ];
	assign fresh_wire_1166[ 12 ] = fresh_wire_2262[ 12 ];
	assign fresh_wire_1166[ 13 ] = fresh_wire_2262[ 13 ];
	assign fresh_wire_1166[ 14 ] = fresh_wire_2262[ 14 ];
	assign fresh_wire_1166[ 15 ] = fresh_wire_2262[ 15 ];
	assign fresh_wire_1168[ 0 ] = fresh_wire_1378[ 0 ];
	assign fresh_wire_1168[ 1 ] = fresh_wire_1378[ 1 ];
	assign fresh_wire_1168[ 2 ] = fresh_wire_1378[ 2 ];
	assign fresh_wire_1168[ 3 ] = fresh_wire_1378[ 3 ];
	assign fresh_wire_1168[ 4 ] = fresh_wire_1378[ 4 ];
	assign fresh_wire_1168[ 5 ] = fresh_wire_1378[ 5 ];
	assign fresh_wire_1168[ 6 ] = fresh_wire_1378[ 6 ];
	assign fresh_wire_1168[ 7 ] = fresh_wire_1378[ 7 ];
	assign fresh_wire_1168[ 8 ] = fresh_wire_1378[ 8 ];
	assign fresh_wire_1168[ 9 ] = fresh_wire_1378[ 9 ];
	assign fresh_wire_1168[ 10 ] = fresh_wire_1378[ 10 ];
	assign fresh_wire_1168[ 11 ] = fresh_wire_1378[ 11 ];
	assign fresh_wire_1168[ 12 ] = fresh_wire_1378[ 12 ];
	assign fresh_wire_1168[ 13 ] = fresh_wire_1378[ 13 ];
	assign fresh_wire_1168[ 14 ] = fresh_wire_1378[ 14 ];
	assign fresh_wire_1168[ 15 ] = fresh_wire_1378[ 15 ];
	assign fresh_wire_1169[ 0 ] = fresh_wire_2263[ 0 ];
	assign fresh_wire_1169[ 1 ] = fresh_wire_2263[ 1 ];
	assign fresh_wire_1169[ 2 ] = fresh_wire_2263[ 2 ];
	assign fresh_wire_1169[ 3 ] = fresh_wire_2263[ 3 ];
	assign fresh_wire_1169[ 4 ] = fresh_wire_2263[ 4 ];
	assign fresh_wire_1169[ 5 ] = fresh_wire_2263[ 5 ];
	assign fresh_wire_1169[ 6 ] = fresh_wire_2263[ 6 ];
	assign fresh_wire_1169[ 7 ] = fresh_wire_2263[ 7 ];
	assign fresh_wire_1169[ 8 ] = fresh_wire_2263[ 8 ];
	assign fresh_wire_1169[ 9 ] = fresh_wire_2263[ 9 ];
	assign fresh_wire_1169[ 10 ] = fresh_wire_2263[ 10 ];
	assign fresh_wire_1169[ 11 ] = fresh_wire_2263[ 11 ];
	assign fresh_wire_1169[ 12 ] = fresh_wire_2263[ 12 ];
	assign fresh_wire_1169[ 13 ] = fresh_wire_2263[ 13 ];
	assign fresh_wire_1169[ 14 ] = fresh_wire_2263[ 14 ];
	assign fresh_wire_1169[ 15 ] = fresh_wire_2263[ 15 ];
	assign fresh_wire_1171[ 0 ] = fresh_wire_1191[ 0 ];
	assign fresh_wire_1172[ 0 ] = fresh_wire_1200[ 0 ];
	assign fresh_wire_1174[ 0 ] = fresh_wire_1348[ 0 ];
	assign fresh_wire_1174[ 1 ] = fresh_wire_1348[ 1 ];
	assign fresh_wire_1175[ 0 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1175[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1177[ 0 ] = fresh_wire_1345[ 0 ];
	assign fresh_wire_1177[ 1 ] = fresh_wire_1345[ 1 ];
	assign fresh_wire_1178[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1178[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1180[ 0 ] = fresh_wire_1638[ 0 ];
	assign fresh_wire_1180[ 1 ] = fresh_wire_1638[ 1 ];
	assign fresh_wire_1181[ 0 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1181[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1183[ 0 ] = fresh_wire_1138[ 0 ];
	assign fresh_wire_1183[ 1 ] = fresh_wire_1138[ 1 ];
	assign fresh_wire_1183[ 2 ] = fresh_wire_1138[ 2 ];
	assign fresh_wire_1183[ 3 ] = fresh_wire_1138[ 3 ];
	assign fresh_wire_1183[ 4 ] = fresh_wire_1138[ 4 ];
	assign fresh_wire_1183[ 5 ] = fresh_wire_1138[ 5 ];
	assign fresh_wire_1183[ 6 ] = fresh_wire_1138[ 6 ];
	assign fresh_wire_1183[ 7 ] = fresh_wire_1138[ 7 ];
	assign fresh_wire_1183[ 8 ] = fresh_wire_1138[ 8 ];
	assign fresh_wire_1183[ 9 ] = fresh_wire_1138[ 9 ];
	assign fresh_wire_1183[ 10 ] = fresh_wire_1138[ 10 ];
	assign fresh_wire_1183[ 11 ] = fresh_wire_1138[ 11 ];
	assign fresh_wire_1183[ 12 ] = fresh_wire_1138[ 12 ];
	assign fresh_wire_1183[ 13 ] = fresh_wire_1138[ 13 ];
	assign fresh_wire_1183[ 14 ] = fresh_wire_1138[ 14 ];
	assign fresh_wire_1183[ 15 ] = fresh_wire_1138[ 15 ];
	assign fresh_wire_1184[ 0 ] = fresh_wire_2264[ 0 ];
	assign fresh_wire_1184[ 1 ] = fresh_wire_2264[ 1 ];
	assign fresh_wire_1184[ 2 ] = fresh_wire_2264[ 2 ];
	assign fresh_wire_1184[ 3 ] = fresh_wire_2264[ 3 ];
	assign fresh_wire_1184[ 4 ] = fresh_wire_2264[ 4 ];
	assign fresh_wire_1184[ 5 ] = fresh_wire_2264[ 5 ];
	assign fresh_wire_1184[ 6 ] = fresh_wire_2264[ 6 ];
	assign fresh_wire_1184[ 7 ] = fresh_wire_2264[ 7 ];
	assign fresh_wire_1184[ 8 ] = fresh_wire_2264[ 8 ];
	assign fresh_wire_1184[ 9 ] = fresh_wire_2264[ 9 ];
	assign fresh_wire_1184[ 10 ] = fresh_wire_2264[ 10 ];
	assign fresh_wire_1184[ 11 ] = fresh_wire_2264[ 11 ];
	assign fresh_wire_1184[ 12 ] = fresh_wire_2264[ 12 ];
	assign fresh_wire_1184[ 13 ] = fresh_wire_2264[ 13 ];
	assign fresh_wire_1184[ 14 ] = fresh_wire_2264[ 14 ];
	assign fresh_wire_1184[ 15 ] = fresh_wire_2264[ 15 ];
	assign fresh_wire_1186[ 0 ] = fresh_wire_1394[ 0 ];
	assign fresh_wire_1187[ 0 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1189[ 0 ] = fresh_wire_1402[ 0 ];
	assign fresh_wire_1190[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1192[ 0 ] = fresh_wire_1650[ 0 ];
	assign fresh_wire_1193[ 0 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1195[ 0 ] = fresh_wire_1258[ 0 ];
	assign fresh_wire_1196[ 0 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1198[ 0 ] = fresh_wire_1374[ 0 ];
	assign fresh_wire_1198[ 1 ] = fresh_wire_1374[ 1 ];
	assign fresh_wire_1199[ 0 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1199[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1201[ 0 ] = fresh_wire_1402[ 0 ];
	assign fresh_wire_1202[ 0 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1204[ 0 ] = fresh_wire_1398[ 0 ];
	assign fresh_wire_1205[ 0 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1207[ 0 ] = fresh_wire_1374[ 0 ];
	assign fresh_wire_1207[ 1 ] = fresh_wire_1374[ 1 ];
	assign fresh_wire_1208[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1208[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1210[ 0 ] = fresh_wire_1335[ 0 ];
	assign fresh_wire_1211[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1213[ 0 ] = fresh_wire_1370[ 0 ];
	assign fresh_wire_1214[ 0 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1216[ 0 ] = fresh_wire_1374[ 0 ];
	assign fresh_wire_1216[ 1 ] = fresh_wire_1374[ 1 ];
	assign fresh_wire_1217[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1217[ 1 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1219[ 0 ] = fresh_wire_1345[ 0 ];
	assign fresh_wire_1219[ 1 ] = fresh_wire_1345[ 1 ];
	assign fresh_wire_1220[ 0 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1220[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1222[ 0 ] = fresh_wire_1170[ 0 ];
	assign fresh_wire_1222[ 1 ] = fresh_wire_1170[ 1 ];
	assign fresh_wire_1222[ 2 ] = fresh_wire_1170[ 2 ];
	assign fresh_wire_1222[ 3 ] = fresh_wire_1170[ 3 ];
	assign fresh_wire_1222[ 4 ] = fresh_wire_1170[ 4 ];
	assign fresh_wire_1222[ 5 ] = fresh_wire_1170[ 5 ];
	assign fresh_wire_1222[ 6 ] = fresh_wire_1170[ 6 ];
	assign fresh_wire_1222[ 7 ] = fresh_wire_1170[ 7 ];
	assign fresh_wire_1222[ 8 ] = fresh_wire_1170[ 8 ];
	assign fresh_wire_1222[ 9 ] = fresh_wire_1170[ 9 ];
	assign fresh_wire_1222[ 10 ] = fresh_wire_1170[ 10 ];
	assign fresh_wire_1222[ 11 ] = fresh_wire_1170[ 11 ];
	assign fresh_wire_1222[ 12 ] = fresh_wire_1170[ 12 ];
	assign fresh_wire_1222[ 13 ] = fresh_wire_1170[ 13 ];
	assign fresh_wire_1222[ 14 ] = fresh_wire_1170[ 14 ];
	assign fresh_wire_1222[ 15 ] = fresh_wire_1170[ 15 ];
	assign fresh_wire_1223[ 0 ] = fresh_wire_2265[ 0 ];
	assign fresh_wire_1223[ 1 ] = fresh_wire_2265[ 1 ];
	assign fresh_wire_1223[ 2 ] = fresh_wire_2265[ 2 ];
	assign fresh_wire_1223[ 3 ] = fresh_wire_2265[ 3 ];
	assign fresh_wire_1223[ 4 ] = fresh_wire_2265[ 4 ];
	assign fresh_wire_1223[ 5 ] = fresh_wire_2265[ 5 ];
	assign fresh_wire_1223[ 6 ] = fresh_wire_2265[ 6 ];
	assign fresh_wire_1223[ 7 ] = fresh_wire_2265[ 7 ];
	assign fresh_wire_1223[ 8 ] = fresh_wire_2265[ 8 ];
	assign fresh_wire_1223[ 9 ] = fresh_wire_2265[ 9 ];
	assign fresh_wire_1223[ 10 ] = fresh_wire_2265[ 10 ];
	assign fresh_wire_1223[ 11 ] = fresh_wire_2265[ 11 ];
	assign fresh_wire_1223[ 12 ] = fresh_wire_2265[ 12 ];
	assign fresh_wire_1223[ 13 ] = fresh_wire_2265[ 13 ];
	assign fresh_wire_1223[ 14 ] = fresh_wire_2265[ 14 ];
	assign fresh_wire_1223[ 15 ] = fresh_wire_2265[ 15 ];
	assign fresh_wire_1225[ 0 ] = fresh_wire_1866[ 0 ];
	assign fresh_wire_1226[ 0 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1228[ 0 ] = fresh_wire_1366[ 0 ];
	assign fresh_wire_1229[ 0 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1231[ 0 ] = fresh_wire_1386[ 0 ];
	assign fresh_wire_1231[ 1 ] = fresh_wire_1386[ 1 ];
	assign fresh_wire_1231[ 2 ] = fresh_wire_1386[ 2 ];
	assign fresh_wire_1231[ 3 ] = fresh_wire_1386[ 3 ];
	assign fresh_wire_1231[ 4 ] = fresh_wire_1386[ 4 ];
	assign fresh_wire_1231[ 5 ] = fresh_wire_1386[ 5 ];
	assign fresh_wire_1231[ 6 ] = fresh_wire_1386[ 6 ];
	assign fresh_wire_1231[ 7 ] = fresh_wire_1386[ 7 ];
	assign fresh_wire_1231[ 8 ] = fresh_wire_1386[ 8 ];
	assign fresh_wire_1231[ 9 ] = fresh_wire_1386[ 9 ];
	assign fresh_wire_1231[ 10 ] = fresh_wire_1386[ 10 ];
	assign fresh_wire_1231[ 11 ] = fresh_wire_1386[ 11 ];
	assign fresh_wire_1231[ 12 ] = fresh_wire_1386[ 12 ];
	assign fresh_wire_1231[ 13 ] = fresh_wire_1386[ 13 ];
	assign fresh_wire_1231[ 14 ] = fresh_wire_1386[ 14 ];
	assign fresh_wire_1231[ 15 ] = fresh_wire_1386[ 15 ];
	assign fresh_wire_1232[ 0 ] = fresh_wire_2267[ 0 ];
	assign fresh_wire_1232[ 1 ] = fresh_wire_2267[ 1 ];
	assign fresh_wire_1232[ 2 ] = fresh_wire_2267[ 2 ];
	assign fresh_wire_1232[ 3 ] = fresh_wire_2267[ 3 ];
	assign fresh_wire_1232[ 4 ] = fresh_wire_2267[ 4 ];
	assign fresh_wire_1232[ 5 ] = fresh_wire_2267[ 5 ];
	assign fresh_wire_1232[ 6 ] = fresh_wire_2267[ 6 ];
	assign fresh_wire_1232[ 7 ] = fresh_wire_2267[ 7 ];
	assign fresh_wire_1232[ 8 ] = fresh_wire_2267[ 8 ];
	assign fresh_wire_1232[ 9 ] = fresh_wire_2267[ 9 ];
	assign fresh_wire_1232[ 10 ] = fresh_wire_2267[ 10 ];
	assign fresh_wire_1232[ 11 ] = fresh_wire_2267[ 11 ];
	assign fresh_wire_1232[ 12 ] = fresh_wire_2267[ 12 ];
	assign fresh_wire_1232[ 13 ] = fresh_wire_2267[ 13 ];
	assign fresh_wire_1232[ 14 ] = fresh_wire_2267[ 14 ];
	assign fresh_wire_1232[ 15 ] = fresh_wire_2267[ 15 ];
	assign fresh_wire_1234[ 0 ] = fresh_wire_1382[ 0 ];
	assign fresh_wire_1234[ 1 ] = fresh_wire_1382[ 1 ];
	assign fresh_wire_1234[ 2 ] = fresh_wire_1382[ 2 ];
	assign fresh_wire_1234[ 3 ] = fresh_wire_1382[ 3 ];
	assign fresh_wire_1234[ 4 ] = fresh_wire_1382[ 4 ];
	assign fresh_wire_1234[ 5 ] = fresh_wire_1382[ 5 ];
	assign fresh_wire_1234[ 6 ] = fresh_wire_1382[ 6 ];
	assign fresh_wire_1234[ 7 ] = fresh_wire_1382[ 7 ];
	assign fresh_wire_1234[ 8 ] = fresh_wire_1382[ 8 ];
	assign fresh_wire_1234[ 9 ] = fresh_wire_1382[ 9 ];
	assign fresh_wire_1234[ 10 ] = fresh_wire_1382[ 10 ];
	assign fresh_wire_1234[ 11 ] = fresh_wire_1382[ 11 ];
	assign fresh_wire_1234[ 12 ] = fresh_wire_1382[ 12 ];
	assign fresh_wire_1234[ 13 ] = fresh_wire_1382[ 13 ];
	assign fresh_wire_1234[ 14 ] = fresh_wire_1382[ 14 ];
	assign fresh_wire_1234[ 15 ] = fresh_wire_1382[ 15 ];
	assign fresh_wire_1235[ 0 ] = fresh_wire_2267[ 0 ];
	assign fresh_wire_1235[ 1 ] = fresh_wire_2267[ 1 ];
	assign fresh_wire_1235[ 2 ] = fresh_wire_2267[ 2 ];
	assign fresh_wire_1235[ 3 ] = fresh_wire_2267[ 3 ];
	assign fresh_wire_1235[ 4 ] = fresh_wire_2267[ 4 ];
	assign fresh_wire_1235[ 5 ] = fresh_wire_2267[ 5 ];
	assign fresh_wire_1235[ 6 ] = fresh_wire_2267[ 6 ];
	assign fresh_wire_1235[ 7 ] = fresh_wire_2267[ 7 ];
	assign fresh_wire_1235[ 8 ] = fresh_wire_2267[ 8 ];
	assign fresh_wire_1235[ 9 ] = fresh_wire_2267[ 9 ];
	assign fresh_wire_1235[ 10 ] = fresh_wire_2267[ 10 ];
	assign fresh_wire_1235[ 11 ] = fresh_wire_2267[ 11 ];
	assign fresh_wire_1235[ 12 ] = fresh_wire_2267[ 12 ];
	assign fresh_wire_1235[ 13 ] = fresh_wire_2267[ 13 ];
	assign fresh_wire_1235[ 14 ] = fresh_wire_2267[ 14 ];
	assign fresh_wire_1235[ 15 ] = fresh_wire_2267[ 15 ];
	assign fresh_wire_1237[ 0 ] = fresh_wire_1167[ 0 ];
	assign fresh_wire_1237[ 1 ] = fresh_wire_1167[ 1 ];
	assign fresh_wire_1237[ 2 ] = fresh_wire_1167[ 2 ];
	assign fresh_wire_1237[ 3 ] = fresh_wire_1167[ 3 ];
	assign fresh_wire_1237[ 4 ] = fresh_wire_1167[ 4 ];
	assign fresh_wire_1237[ 5 ] = fresh_wire_1167[ 5 ];
	assign fresh_wire_1237[ 6 ] = fresh_wire_1167[ 6 ];
	assign fresh_wire_1237[ 7 ] = fresh_wire_1167[ 7 ];
	assign fresh_wire_1237[ 8 ] = fresh_wire_1167[ 8 ];
	assign fresh_wire_1237[ 9 ] = fresh_wire_1167[ 9 ];
	assign fresh_wire_1237[ 10 ] = fresh_wire_1167[ 10 ];
	assign fresh_wire_1237[ 11 ] = fresh_wire_1167[ 11 ];
	assign fresh_wire_1237[ 12 ] = fresh_wire_1167[ 12 ];
	assign fresh_wire_1237[ 13 ] = fresh_wire_1167[ 13 ];
	assign fresh_wire_1237[ 14 ] = fresh_wire_1167[ 14 ];
	assign fresh_wire_1237[ 15 ] = fresh_wire_1167[ 15 ];
	assign fresh_wire_1238[ 0 ] = fresh_wire_2266[ 0 ];
	assign fresh_wire_1238[ 1 ] = fresh_wire_2266[ 1 ];
	assign fresh_wire_1238[ 2 ] = fresh_wire_2266[ 2 ];
	assign fresh_wire_1238[ 3 ] = fresh_wire_2266[ 3 ];
	assign fresh_wire_1238[ 4 ] = fresh_wire_2266[ 4 ];
	assign fresh_wire_1238[ 5 ] = fresh_wire_2266[ 5 ];
	assign fresh_wire_1238[ 6 ] = fresh_wire_2266[ 6 ];
	assign fresh_wire_1238[ 7 ] = fresh_wire_2266[ 7 ];
	assign fresh_wire_1238[ 8 ] = fresh_wire_2266[ 8 ];
	assign fresh_wire_1238[ 9 ] = fresh_wire_2266[ 9 ];
	assign fresh_wire_1238[ 10 ] = fresh_wire_2266[ 10 ];
	assign fresh_wire_1238[ 11 ] = fresh_wire_2266[ 11 ];
	assign fresh_wire_1238[ 12 ] = fresh_wire_2266[ 12 ];
	assign fresh_wire_1238[ 13 ] = fresh_wire_2266[ 13 ];
	assign fresh_wire_1238[ 14 ] = fresh_wire_2266[ 14 ];
	assign fresh_wire_1238[ 15 ] = fresh_wire_2266[ 15 ];
	assign fresh_wire_1240[ 0 ] = fresh_wire_1176[ 0 ];
	assign fresh_wire_1242[ 0 ] = fresh_wire_1241[ 0 ];
	assign fresh_wire_1243[ 0 ] = fresh_wire_1246[ 0 ];
	assign fresh_wire_1245[ 0 ] = fresh_wire_1179[ 0 ];
	assign fresh_wire_1247[ 0 ] = fresh_wire_1244[ 0 ];
	assign fresh_wire_1249[ 0 ] = fresh_wire_1248[ 0 ];
	assign fresh_wire_1250[ 0 ] = fresh_wire_1253[ 0 ];
	assign fresh_wire_1252[ 0 ] = fresh_wire_1182[ 0 ];
	assign fresh_wire_1254[ 0 ] = fresh_wire_1251[ 0 ];
	assign fresh_wire_1256[ 0 ] = fresh_wire_1255[ 0 ];
	assign fresh_wire_1257[ 0 ] = fresh_wire_1260[ 0 ];
	assign fresh_wire_1259[ 0 ] = fresh_wire_1185[ 0 ];
	assign fresh_wire_1261[ 0 ] = fresh_wire_1209[ 0 ];
	assign fresh_wire_1263[ 0 ] = fresh_wire_1262[ 0 ];
	assign fresh_wire_1264[ 0 ] = fresh_wire_2314[ 0 ];
	assign fresh_wire_1266[ 0 ] = fresh_wire_1265[ 0 ];
	assign fresh_wire_1268[ 0 ] = fresh_wire_1267[ 0 ];
	assign fresh_wire_1269[ 0 ] = fresh_wire_1272[ 0 ];
	assign fresh_wire_1271[ 0 ] = fresh_wire_1212[ 0 ];
	assign fresh_wire_1273[ 0 ] = fresh_wire_1200[ 0 ];
	assign fresh_wire_1275[ 0 ] = fresh_wire_1274[ 0 ];
	assign fresh_wire_1276[ 0 ] = fresh_wire_2315[ 0 ];
	assign fresh_wire_1278[ 0 ] = fresh_wire_1277[ 0 ];
	assign fresh_wire_1280[ 0 ] = fresh_wire_1279[ 0 ];
	assign fresh_wire_1281[ 0 ] = fresh_wire_1284[ 0 ];
	assign fresh_wire_1283[ 0 ] = fresh_wire_1338[ 0 ];
	assign fresh_wire_1285[ 0 ] = fresh_wire_1200[ 0 ];
	assign fresh_wire_1287[ 0 ] = fresh_wire_1286[ 0 ];
	assign fresh_wire_1288[ 0 ] = fresh_wire_1291[ 0 ];
	assign fresh_wire_1290[ 0 ] = fresh_wire_1239[ 0 ];
	assign fresh_wire_1292[ 0 ] = fresh_wire_2316[ 0 ];
	assign fresh_wire_1293[ 0 ] = fresh_wire_1296[ 0 ];
	assign fresh_wire_1295[ 0 ] = fresh_wire_1212[ 0 ];
	assign fresh_wire_1297[ 0 ] = fresh_wire_1218[ 0 ];
	assign fresh_wire_1299[ 0 ] = fresh_wire_1298[ 0 ];
	assign fresh_wire_1300[ 0 ] = fresh_wire_2317[ 0 ];
	assign fresh_wire_1302[ 0 ] = fresh_wire_1176[ 0 ];
	assign fresh_wire_1304[ 0 ] = fresh_wire_1303[ 0 ];
	assign fresh_wire_1305[ 0 ] = fresh_wire_1308[ 0 ];
	assign fresh_wire_1307[ 0 ] = fresh_wire_1179[ 0 ];
	assign fresh_wire_1309[ 0 ] = fresh_wire_1306[ 0 ];
	assign fresh_wire_1311[ 0 ] = fresh_wire_1310[ 0 ];
	assign fresh_wire_1312[ 0 ] = fresh_wire_1315[ 0 ];
	assign fresh_wire_1314[ 0 ] = fresh_wire_1182[ 0 ];
	assign fresh_wire_1316[ 0 ] = fresh_wire_1313[ 0 ];
	assign fresh_wire_1318[ 0 ] = fresh_wire_1317[ 0 ];
	assign fresh_wire_1319[ 0 ] = fresh_wire_1322[ 0 ];
	assign fresh_wire_1321[ 0 ] = fresh_wire_1224[ 0 ];
	assign fresh_wire_1323[ 0 ] = fresh_wire_1227[ 0 ];
	assign fresh_wire_1325[ 0 ] = fresh_wire_1324[ 0 ];
	assign fresh_wire_1326[ 0 ] = fresh_wire_2318[ 0 ];
	assign fresh_wire_1328[ 0 ] = fresh_wire_1335[ 0 ];
	assign fresh_wire_1330[ 0 ] = fresh_wire_2319[ 0 ];
	assign fresh_wire_1331[ 0 ] = fresh_wire_1329[ 0 ];
	assign fresh_wire_1333[ 0 ] = fresh_wire_1143[ 0 ];
	assign fresh_wire_1333[ 1 ] = fresh_wire_1143[ 1 ];
	assign fresh_wire_1333[ 2 ] = fresh_wire_1143[ 2 ];
	assign fresh_wire_1333[ 3 ] = fresh_wire_1143[ 3 ];
	assign fresh_wire_1333[ 4 ] = fresh_wire_1143[ 4 ];
	assign fresh_wire_1333[ 5 ] = fresh_wire_1143[ 5 ];
	assign fresh_wire_1333[ 6 ] = fresh_wire_1143[ 6 ];
	assign fresh_wire_1333[ 7 ] = fresh_wire_1143[ 7 ];
	assign fresh_wire_1333[ 8 ] = fresh_wire_1143[ 8 ];
	assign fresh_wire_1333[ 9 ] = fresh_wire_1143[ 9 ];
	assign fresh_wire_1333[ 10 ] = fresh_wire_1143[ 10 ];
	assign fresh_wire_1333[ 11 ] = fresh_wire_1143[ 11 ];
	assign fresh_wire_1333[ 12 ] = fresh_wire_1143[ 12 ];
	assign fresh_wire_1333[ 13 ] = fresh_wire_1143[ 13 ];
	assign fresh_wire_1333[ 14 ] = fresh_wire_1143[ 14 ];
	assign fresh_wire_1333[ 15 ] = fresh_wire_1143[ 15 ];
	assign fresh_wire_1334[ 0 ] = fresh_wire_2268[ 0 ];
	assign fresh_wire_1334[ 1 ] = fresh_wire_2268[ 1 ];
	assign fresh_wire_1334[ 2 ] = fresh_wire_2268[ 2 ];
	assign fresh_wire_1334[ 3 ] = fresh_wire_2268[ 3 ];
	assign fresh_wire_1334[ 4 ] = fresh_wire_2268[ 4 ];
	assign fresh_wire_1334[ 5 ] = fresh_wire_2268[ 5 ];
	assign fresh_wire_1334[ 6 ] = fresh_wire_2268[ 6 ];
	assign fresh_wire_1334[ 7 ] = fresh_wire_2268[ 7 ];
	assign fresh_wire_1334[ 8 ] = fresh_wire_2268[ 8 ];
	assign fresh_wire_1334[ 9 ] = fresh_wire_2268[ 9 ];
	assign fresh_wire_1334[ 10 ] = fresh_wire_2268[ 10 ];
	assign fresh_wire_1334[ 11 ] = fresh_wire_2268[ 11 ];
	assign fresh_wire_1334[ 12 ] = fresh_wire_2268[ 12 ];
	assign fresh_wire_1334[ 13 ] = fresh_wire_2268[ 13 ];
	assign fresh_wire_1334[ 14 ] = fresh_wire_2268[ 14 ];
	assign fresh_wire_1334[ 15 ] = fresh_wire_2268[ 15 ];
	assign fresh_wire_1336[ 0 ] = fresh_wire_1161[ 0 ];
	assign fresh_wire_1336[ 1 ] = fresh_wire_1161[ 1 ];
	assign fresh_wire_1336[ 2 ] = fresh_wire_1161[ 2 ];
	assign fresh_wire_1336[ 3 ] = fresh_wire_1161[ 3 ];
	assign fresh_wire_1336[ 4 ] = fresh_wire_1161[ 4 ];
	assign fresh_wire_1336[ 5 ] = fresh_wire_1161[ 5 ];
	assign fresh_wire_1336[ 6 ] = fresh_wire_1161[ 6 ];
	assign fresh_wire_1336[ 7 ] = fresh_wire_1161[ 7 ];
	assign fresh_wire_1336[ 8 ] = fresh_wire_1161[ 8 ];
	assign fresh_wire_1336[ 9 ] = fresh_wire_1161[ 9 ];
	assign fresh_wire_1336[ 10 ] = fresh_wire_1161[ 10 ];
	assign fresh_wire_1336[ 11 ] = fresh_wire_1161[ 11 ];
	assign fresh_wire_1336[ 12 ] = fresh_wire_1161[ 12 ];
	assign fresh_wire_1336[ 13 ] = fresh_wire_1161[ 13 ];
	assign fresh_wire_1336[ 14 ] = fresh_wire_1161[ 14 ];
	assign fresh_wire_1336[ 15 ] = fresh_wire_1161[ 15 ];
	assign fresh_wire_1337[ 0 ] = fresh_wire_2266[ 0 ];
	assign fresh_wire_1337[ 1 ] = fresh_wire_2266[ 1 ];
	assign fresh_wire_1337[ 2 ] = fresh_wire_2266[ 2 ];
	assign fresh_wire_1337[ 3 ] = fresh_wire_2266[ 3 ];
	assign fresh_wire_1337[ 4 ] = fresh_wire_2266[ 4 ];
	assign fresh_wire_1337[ 5 ] = fresh_wire_2266[ 5 ];
	assign fresh_wire_1337[ 6 ] = fresh_wire_2266[ 6 ];
	assign fresh_wire_1337[ 7 ] = fresh_wire_2266[ 7 ];
	assign fresh_wire_1337[ 8 ] = fresh_wire_2266[ 8 ];
	assign fresh_wire_1337[ 9 ] = fresh_wire_2266[ 9 ];
	assign fresh_wire_1337[ 10 ] = fresh_wire_2266[ 10 ];
	assign fresh_wire_1337[ 11 ] = fresh_wire_2266[ 11 ];
	assign fresh_wire_1337[ 12 ] = fresh_wire_2266[ 12 ];
	assign fresh_wire_1337[ 13 ] = fresh_wire_2266[ 13 ];
	assign fresh_wire_1337[ 14 ] = fresh_wire_2266[ 14 ];
	assign fresh_wire_1337[ 15 ] = fresh_wire_2266[ 15 ];
	assign fresh_wire_1339[ 0 ] = fresh_wire_1402[ 0 ];
	assign fresh_wire_1341[ 0 ] = fresh_wire_1332[ 0 ];
	assign fresh_wire_1343[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1344[ 0 ] = fresh_wire_1374[ 0 ];
	assign fresh_wire_1344[ 1 ] = fresh_wire_1374[ 1 ];
	assign fresh_wire_1346[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1347[ 0 ] = fresh_wire_1345[ 0 ];
	assign fresh_wire_1347[ 1 ] = fresh_wire_1345[ 1 ];
	assign fresh_wire_1349[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1350[ 0 ] = fresh_wire_1850[ 0 ];
	assign fresh_wire_1350[ 1 ] = fresh_wire_1850[ 1 ];
	assign fresh_wire_1350[ 2 ] = fresh_wire_1850[ 2 ];
	assign fresh_wire_1350[ 3 ] = fresh_wire_1850[ 3 ];
	assign fresh_wire_1350[ 4 ] = fresh_wire_1850[ 4 ];
	assign fresh_wire_1350[ 5 ] = fresh_wire_1850[ 5 ];
	assign fresh_wire_1350[ 6 ] = fresh_wire_1850[ 6 ];
	assign fresh_wire_1350[ 7 ] = fresh_wire_1850[ 7 ];
	assign fresh_wire_1350[ 8 ] = fresh_wire_1850[ 8 ];
	assign fresh_wire_1350[ 9 ] = fresh_wire_1850[ 9 ];
	assign fresh_wire_1350[ 10 ] = fresh_wire_1850[ 10 ];
	assign fresh_wire_1350[ 11 ] = fresh_wire_1850[ 11 ];
	assign fresh_wire_1350[ 12 ] = fresh_wire_1850[ 12 ];
	assign fresh_wire_1350[ 13 ] = fresh_wire_1850[ 13 ];
	assign fresh_wire_1350[ 14 ] = fresh_wire_1850[ 14 ];
	assign fresh_wire_1350[ 15 ] = fresh_wire_1850[ 15 ];
	assign fresh_wire_1352[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1353[ 0 ] = fresh_wire_1427[ 0 ];
	assign fresh_wire_1355[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1356[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_1357[ 0 ] = fresh_wire_1423[ 0 ];
	assign fresh_wire_1359[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1360[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_1361[ 0 ] = fresh_wire_1415[ 0 ];
	assign fresh_wire_1363[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1364[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_1365[ 0 ] = fresh_wire_1507[ 0 ];
	assign fresh_wire_1367[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1368[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_1369[ 0 ] = fresh_wire_1483[ 0 ];
	assign fresh_wire_1371[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1372[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_1373[ 0 ] = fresh_wire_1467[ 0 ];
	assign fresh_wire_1373[ 1 ] = fresh_wire_1467[ 1 ];
	assign fresh_wire_1375[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1376[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_1377[ 0 ] = fresh_wire_1443[ 0 ];
	assign fresh_wire_1377[ 1 ] = fresh_wire_1443[ 1 ];
	assign fresh_wire_1377[ 2 ] = fresh_wire_1443[ 2 ];
	assign fresh_wire_1377[ 3 ] = fresh_wire_1443[ 3 ];
	assign fresh_wire_1377[ 4 ] = fresh_wire_1443[ 4 ];
	assign fresh_wire_1377[ 5 ] = fresh_wire_1443[ 5 ];
	assign fresh_wire_1377[ 6 ] = fresh_wire_1443[ 6 ];
	assign fresh_wire_1377[ 7 ] = fresh_wire_1443[ 7 ];
	assign fresh_wire_1377[ 8 ] = fresh_wire_1443[ 8 ];
	assign fresh_wire_1377[ 9 ] = fresh_wire_1443[ 9 ];
	assign fresh_wire_1377[ 10 ] = fresh_wire_1443[ 10 ];
	assign fresh_wire_1377[ 11 ] = fresh_wire_1443[ 11 ];
	assign fresh_wire_1377[ 12 ] = fresh_wire_1443[ 12 ];
	assign fresh_wire_1377[ 13 ] = fresh_wire_1443[ 13 ];
	assign fresh_wire_1377[ 14 ] = fresh_wire_1443[ 14 ];
	assign fresh_wire_1377[ 15 ] = fresh_wire_1443[ 15 ];
	assign fresh_wire_1379[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1380[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_1381[ 0 ] = fresh_wire_1543[ 0 ];
	assign fresh_wire_1381[ 1 ] = fresh_wire_1543[ 1 ];
	assign fresh_wire_1381[ 2 ] = fresh_wire_1543[ 2 ];
	assign fresh_wire_1381[ 3 ] = fresh_wire_1543[ 3 ];
	assign fresh_wire_1381[ 4 ] = fresh_wire_1543[ 4 ];
	assign fresh_wire_1381[ 5 ] = fresh_wire_1543[ 5 ];
	assign fresh_wire_1381[ 6 ] = fresh_wire_1543[ 6 ];
	assign fresh_wire_1381[ 7 ] = fresh_wire_1543[ 7 ];
	assign fresh_wire_1381[ 8 ] = fresh_wire_1543[ 8 ];
	assign fresh_wire_1381[ 9 ] = fresh_wire_1543[ 9 ];
	assign fresh_wire_1381[ 10 ] = fresh_wire_1543[ 10 ];
	assign fresh_wire_1381[ 11 ] = fresh_wire_1543[ 11 ];
	assign fresh_wire_1381[ 12 ] = fresh_wire_1543[ 12 ];
	assign fresh_wire_1381[ 13 ] = fresh_wire_1543[ 13 ];
	assign fresh_wire_1381[ 14 ] = fresh_wire_1543[ 14 ];
	assign fresh_wire_1381[ 15 ] = fresh_wire_1543[ 15 ];
	assign fresh_wire_1383[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1384[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_1385[ 0 ] = fresh_wire_1531[ 0 ];
	assign fresh_wire_1385[ 1 ] = fresh_wire_1531[ 1 ];
	assign fresh_wire_1385[ 2 ] = fresh_wire_1531[ 2 ];
	assign fresh_wire_1385[ 3 ] = fresh_wire_1531[ 3 ];
	assign fresh_wire_1385[ 4 ] = fresh_wire_1531[ 4 ];
	assign fresh_wire_1385[ 5 ] = fresh_wire_1531[ 5 ];
	assign fresh_wire_1385[ 6 ] = fresh_wire_1531[ 6 ];
	assign fresh_wire_1385[ 7 ] = fresh_wire_1531[ 7 ];
	assign fresh_wire_1385[ 8 ] = fresh_wire_1531[ 8 ];
	assign fresh_wire_1385[ 9 ] = fresh_wire_1531[ 9 ];
	assign fresh_wire_1385[ 10 ] = fresh_wire_1531[ 10 ];
	assign fresh_wire_1385[ 11 ] = fresh_wire_1531[ 11 ];
	assign fresh_wire_1385[ 12 ] = fresh_wire_1531[ 12 ];
	assign fresh_wire_1385[ 13 ] = fresh_wire_1531[ 13 ];
	assign fresh_wire_1385[ 14 ] = fresh_wire_1531[ 14 ];
	assign fresh_wire_1385[ 15 ] = fresh_wire_1531[ 15 ];
	assign fresh_wire_1387[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1388[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_1389[ 0 ] = fresh_wire_1519[ 0 ];
	assign fresh_wire_1389[ 1 ] = fresh_wire_1519[ 1 ];
	assign fresh_wire_1389[ 2 ] = fresh_wire_1519[ 2 ];
	assign fresh_wire_1389[ 3 ] = fresh_wire_1519[ 3 ];
	assign fresh_wire_1389[ 4 ] = fresh_wire_1519[ 4 ];
	assign fresh_wire_1389[ 5 ] = fresh_wire_1519[ 5 ];
	assign fresh_wire_1389[ 6 ] = fresh_wire_1519[ 6 ];
	assign fresh_wire_1389[ 7 ] = fresh_wire_1519[ 7 ];
	assign fresh_wire_1389[ 8 ] = fresh_wire_1519[ 8 ];
	assign fresh_wire_1389[ 9 ] = fresh_wire_1519[ 9 ];
	assign fresh_wire_1389[ 10 ] = fresh_wire_1519[ 10 ];
	assign fresh_wire_1389[ 11 ] = fresh_wire_1519[ 11 ];
	assign fresh_wire_1389[ 12 ] = fresh_wire_1519[ 12 ];
	assign fresh_wire_1389[ 13 ] = fresh_wire_1519[ 13 ];
	assign fresh_wire_1389[ 14 ] = fresh_wire_1519[ 14 ];
	assign fresh_wire_1389[ 15 ] = fresh_wire_1519[ 15 ];
	assign fresh_wire_1391[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1392[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_1393[ 0 ] = fresh_wire_1563[ 0 ];
	assign fresh_wire_1395[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1396[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_1397[ 0 ] = fresh_wire_1551[ 0 ];
	assign fresh_wire_1399[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1400[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_1401[ 0 ] = fresh_wire_1340[ 0 ];
	assign fresh_wire_1403[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1404[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_1405[ 0 ] = fresh_wire_1386[ 0 ];
	assign fresh_wire_1405[ 1 ] = fresh_wire_1386[ 1 ];
	assign fresh_wire_1405[ 2 ] = fresh_wire_1386[ 2 ];
	assign fresh_wire_1405[ 3 ] = fresh_wire_1386[ 3 ];
	assign fresh_wire_1405[ 4 ] = fresh_wire_1386[ 4 ];
	assign fresh_wire_1405[ 5 ] = fresh_wire_1386[ 5 ];
	assign fresh_wire_1405[ 6 ] = fresh_wire_1386[ 6 ];
	assign fresh_wire_1405[ 7 ] = fresh_wire_1386[ 7 ];
	assign fresh_wire_1405[ 8 ] = fresh_wire_1386[ 8 ];
	assign fresh_wire_1405[ 9 ] = fresh_wire_1386[ 9 ];
	assign fresh_wire_1405[ 10 ] = fresh_wire_1386[ 10 ];
	assign fresh_wire_1405[ 11 ] = fresh_wire_1386[ 11 ];
	assign fresh_wire_1405[ 12 ] = fresh_wire_1386[ 12 ];
	assign fresh_wire_1405[ 13 ] = fresh_wire_1386[ 13 ];
	assign fresh_wire_1405[ 14 ] = fresh_wire_1386[ 14 ];
	assign fresh_wire_1405[ 15 ] = fresh_wire_1386[ 15 ];
	assign fresh_wire_1406[ 0 ] = fresh_wire_1382[ 0 ];
	assign fresh_wire_1406[ 1 ] = fresh_wire_1382[ 1 ];
	assign fresh_wire_1406[ 2 ] = fresh_wire_1382[ 2 ];
	assign fresh_wire_1406[ 3 ] = fresh_wire_1382[ 3 ];
	assign fresh_wire_1406[ 4 ] = fresh_wire_1382[ 4 ];
	assign fresh_wire_1406[ 5 ] = fresh_wire_1382[ 5 ];
	assign fresh_wire_1406[ 6 ] = fresh_wire_1382[ 6 ];
	assign fresh_wire_1406[ 7 ] = fresh_wire_1382[ 7 ];
	assign fresh_wire_1406[ 8 ] = fresh_wire_1382[ 8 ];
	assign fresh_wire_1406[ 9 ] = fresh_wire_1382[ 9 ];
	assign fresh_wire_1406[ 10 ] = fresh_wire_1382[ 10 ];
	assign fresh_wire_1406[ 11 ] = fresh_wire_1382[ 11 ];
	assign fresh_wire_1406[ 12 ] = fresh_wire_1382[ 12 ];
	assign fresh_wire_1406[ 13 ] = fresh_wire_1382[ 13 ];
	assign fresh_wire_1406[ 14 ] = fresh_wire_1382[ 14 ];
	assign fresh_wire_1406[ 15 ] = fresh_wire_1382[ 15 ];
	assign fresh_wire_1408[ 0 ] = fresh_wire_1191[ 0 ];
	assign fresh_wire_1409[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1410[ 0 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1412[ 0 ] = fresh_wire_1221[ 0 ];
	assign fresh_wire_1413[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1414[ 0 ] = fresh_wire_1411[ 0 ];
	assign fresh_wire_1416[ 0 ] = fresh_wire_1191[ 0 ];
	assign fresh_wire_1417[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1418[ 0 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1420[ 0 ] = fresh_wire_1320[ 0 ];
	assign fresh_wire_1421[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1422[ 0 ] = fresh_wire_1419[ 0 ];
	assign fresh_wire_1424[ 0 ] = fresh_wire_1191[ 0 ];
	assign fresh_wire_1425[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1426[ 0 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1428[ 0 ] = fresh_wire_1327[ 0 ];
	assign fresh_wire_1429[ 0 ] = fresh_wire_1378[ 0 ];
	assign fresh_wire_1429[ 1 ] = fresh_wire_1378[ 1 ];
	assign fresh_wire_1429[ 2 ] = fresh_wire_1378[ 2 ];
	assign fresh_wire_1429[ 3 ] = fresh_wire_1378[ 3 ];
	assign fresh_wire_1429[ 4 ] = fresh_wire_1378[ 4 ];
	assign fresh_wire_1429[ 5 ] = fresh_wire_1378[ 5 ];
	assign fresh_wire_1429[ 6 ] = fresh_wire_1378[ 6 ];
	assign fresh_wire_1429[ 7 ] = fresh_wire_1378[ 7 ];
	assign fresh_wire_1429[ 8 ] = fresh_wire_1378[ 8 ];
	assign fresh_wire_1429[ 9 ] = fresh_wire_1378[ 9 ];
	assign fresh_wire_1429[ 10 ] = fresh_wire_1378[ 10 ];
	assign fresh_wire_1429[ 11 ] = fresh_wire_1378[ 11 ];
	assign fresh_wire_1429[ 12 ] = fresh_wire_1378[ 12 ];
	assign fresh_wire_1429[ 13 ] = fresh_wire_1378[ 13 ];
	assign fresh_wire_1429[ 14 ] = fresh_wire_1378[ 14 ];
	assign fresh_wire_1429[ 15 ] = fresh_wire_1378[ 15 ];
	assign fresh_wire_1430[ 0 ] = fresh_wire_1164[ 0 ];
	assign fresh_wire_1430[ 1 ] = fresh_wire_1164[ 1 ];
	assign fresh_wire_1430[ 2 ] = fresh_wire_1164[ 2 ];
	assign fresh_wire_1430[ 3 ] = fresh_wire_1164[ 3 ];
	assign fresh_wire_1430[ 4 ] = fresh_wire_1164[ 4 ];
	assign fresh_wire_1430[ 5 ] = fresh_wire_1164[ 5 ];
	assign fresh_wire_1430[ 6 ] = fresh_wire_1164[ 6 ];
	assign fresh_wire_1430[ 7 ] = fresh_wire_1164[ 7 ];
	assign fresh_wire_1430[ 8 ] = fresh_wire_1164[ 8 ];
	assign fresh_wire_1430[ 9 ] = fresh_wire_1164[ 9 ];
	assign fresh_wire_1430[ 10 ] = fresh_wire_1164[ 10 ];
	assign fresh_wire_1430[ 11 ] = fresh_wire_1164[ 11 ];
	assign fresh_wire_1430[ 12 ] = fresh_wire_1164[ 12 ];
	assign fresh_wire_1430[ 13 ] = fresh_wire_1164[ 13 ];
	assign fresh_wire_1430[ 14 ] = fresh_wire_1164[ 14 ];
	assign fresh_wire_1430[ 15 ] = fresh_wire_1164[ 15 ];
	assign fresh_wire_1432[ 0 ] = fresh_wire_1289[ 0 ];
	assign fresh_wire_1433[ 0 ] = fresh_wire_1431[ 0 ];
	assign fresh_wire_1433[ 1 ] = fresh_wire_1431[ 1 ];
	assign fresh_wire_1433[ 2 ] = fresh_wire_1431[ 2 ];
	assign fresh_wire_1433[ 3 ] = fresh_wire_1431[ 3 ];
	assign fresh_wire_1433[ 4 ] = fresh_wire_1431[ 4 ];
	assign fresh_wire_1433[ 5 ] = fresh_wire_1431[ 5 ];
	assign fresh_wire_1433[ 6 ] = fresh_wire_1431[ 6 ];
	assign fresh_wire_1433[ 7 ] = fresh_wire_1431[ 7 ];
	assign fresh_wire_1433[ 8 ] = fresh_wire_1431[ 8 ];
	assign fresh_wire_1433[ 9 ] = fresh_wire_1431[ 9 ];
	assign fresh_wire_1433[ 10 ] = fresh_wire_1431[ 10 ];
	assign fresh_wire_1433[ 11 ] = fresh_wire_1431[ 11 ];
	assign fresh_wire_1433[ 12 ] = fresh_wire_1431[ 12 ];
	assign fresh_wire_1433[ 13 ] = fresh_wire_1431[ 13 ];
	assign fresh_wire_1433[ 14 ] = fresh_wire_1431[ 14 ];
	assign fresh_wire_1433[ 15 ] = fresh_wire_1431[ 15 ];
	assign fresh_wire_1434[ 0 ] = fresh_wire_1576[ 0 ];
	assign fresh_wire_1434[ 1 ] = fresh_wire_1576[ 1 ];
	assign fresh_wire_1434[ 2 ] = fresh_wire_1576[ 2 ];
	assign fresh_wire_1434[ 3 ] = fresh_wire_1576[ 3 ];
	assign fresh_wire_1434[ 4 ] = fresh_wire_1576[ 4 ];
	assign fresh_wire_1434[ 5 ] = fresh_wire_1576[ 5 ];
	assign fresh_wire_1434[ 6 ] = fresh_wire_1576[ 6 ];
	assign fresh_wire_1434[ 7 ] = fresh_wire_1576[ 7 ];
	assign fresh_wire_1434[ 8 ] = fresh_wire_1576[ 8 ];
	assign fresh_wire_1434[ 9 ] = fresh_wire_1576[ 9 ];
	assign fresh_wire_1434[ 10 ] = fresh_wire_1576[ 10 ];
	assign fresh_wire_1434[ 11 ] = fresh_wire_1576[ 11 ];
	assign fresh_wire_1434[ 12 ] = fresh_wire_1576[ 12 ];
	assign fresh_wire_1434[ 13 ] = fresh_wire_1576[ 13 ];
	assign fresh_wire_1434[ 14 ] = fresh_wire_1576[ 14 ];
	assign fresh_wire_1434[ 15 ] = fresh_wire_1576[ 15 ];
	assign fresh_wire_1436[ 0 ] = fresh_wire_1282[ 0 ];
	assign fresh_wire_1437[ 0 ] = fresh_wire_1435[ 0 ];
	assign fresh_wire_1437[ 1 ] = fresh_wire_1435[ 1 ];
	assign fresh_wire_1437[ 2 ] = fresh_wire_1435[ 2 ];
	assign fresh_wire_1437[ 3 ] = fresh_wire_1435[ 3 ];
	assign fresh_wire_1437[ 4 ] = fresh_wire_1435[ 4 ];
	assign fresh_wire_1437[ 5 ] = fresh_wire_1435[ 5 ];
	assign fresh_wire_1437[ 6 ] = fresh_wire_1435[ 6 ];
	assign fresh_wire_1437[ 7 ] = fresh_wire_1435[ 7 ];
	assign fresh_wire_1437[ 8 ] = fresh_wire_1435[ 8 ];
	assign fresh_wire_1437[ 9 ] = fresh_wire_1435[ 9 ];
	assign fresh_wire_1437[ 10 ] = fresh_wire_1435[ 10 ];
	assign fresh_wire_1437[ 11 ] = fresh_wire_1435[ 11 ];
	assign fresh_wire_1437[ 12 ] = fresh_wire_1435[ 12 ];
	assign fresh_wire_1437[ 13 ] = fresh_wire_1435[ 13 ];
	assign fresh_wire_1437[ 14 ] = fresh_wire_1435[ 14 ];
	assign fresh_wire_1437[ 15 ] = fresh_wire_1435[ 15 ];
	assign fresh_wire_1438[ 0 ] = fresh_wire_1378[ 0 ];
	assign fresh_wire_1438[ 1 ] = fresh_wire_1378[ 1 ];
	assign fresh_wire_1438[ 2 ] = fresh_wire_1378[ 2 ];
	assign fresh_wire_1438[ 3 ] = fresh_wire_1378[ 3 ];
	assign fresh_wire_1438[ 4 ] = fresh_wire_1378[ 4 ];
	assign fresh_wire_1438[ 5 ] = fresh_wire_1378[ 5 ];
	assign fresh_wire_1438[ 6 ] = fresh_wire_1378[ 6 ];
	assign fresh_wire_1438[ 7 ] = fresh_wire_1378[ 7 ];
	assign fresh_wire_1438[ 8 ] = fresh_wire_1378[ 8 ];
	assign fresh_wire_1438[ 9 ] = fresh_wire_1378[ 9 ];
	assign fresh_wire_1438[ 10 ] = fresh_wire_1378[ 10 ];
	assign fresh_wire_1438[ 11 ] = fresh_wire_1378[ 11 ];
	assign fresh_wire_1438[ 12 ] = fresh_wire_1378[ 12 ];
	assign fresh_wire_1438[ 13 ] = fresh_wire_1378[ 13 ];
	assign fresh_wire_1438[ 14 ] = fresh_wire_1378[ 14 ];
	assign fresh_wire_1438[ 15 ] = fresh_wire_1378[ 15 ];
	assign fresh_wire_1440[ 0 ] = fresh_wire_1270[ 0 ];
	assign fresh_wire_1441[ 0 ] = fresh_wire_1378[ 0 ];
	assign fresh_wire_1441[ 1 ] = fresh_wire_1378[ 1 ];
	assign fresh_wire_1441[ 2 ] = fresh_wire_1378[ 2 ];
	assign fresh_wire_1441[ 3 ] = fresh_wire_1378[ 3 ];
	assign fresh_wire_1441[ 4 ] = fresh_wire_1378[ 4 ];
	assign fresh_wire_1441[ 5 ] = fresh_wire_1378[ 5 ];
	assign fresh_wire_1441[ 6 ] = fresh_wire_1378[ 6 ];
	assign fresh_wire_1441[ 7 ] = fresh_wire_1378[ 7 ];
	assign fresh_wire_1441[ 8 ] = fresh_wire_1378[ 8 ];
	assign fresh_wire_1441[ 9 ] = fresh_wire_1378[ 9 ];
	assign fresh_wire_1441[ 10 ] = fresh_wire_1378[ 10 ];
	assign fresh_wire_1441[ 11 ] = fresh_wire_1378[ 11 ];
	assign fresh_wire_1441[ 12 ] = fresh_wire_1378[ 12 ];
	assign fresh_wire_1441[ 13 ] = fresh_wire_1378[ 13 ];
	assign fresh_wire_1441[ 14 ] = fresh_wire_1378[ 14 ];
	assign fresh_wire_1441[ 15 ] = fresh_wire_1378[ 15 ];
	assign fresh_wire_1442[ 0 ] = fresh_wire_1439[ 0 ];
	assign fresh_wire_1442[ 1 ] = fresh_wire_1439[ 1 ];
	assign fresh_wire_1442[ 2 ] = fresh_wire_1439[ 2 ];
	assign fresh_wire_1442[ 3 ] = fresh_wire_1439[ 3 ];
	assign fresh_wire_1442[ 4 ] = fresh_wire_1439[ 4 ];
	assign fresh_wire_1442[ 5 ] = fresh_wire_1439[ 5 ];
	assign fresh_wire_1442[ 6 ] = fresh_wire_1439[ 6 ];
	assign fresh_wire_1442[ 7 ] = fresh_wire_1439[ 7 ];
	assign fresh_wire_1442[ 8 ] = fresh_wire_1439[ 8 ];
	assign fresh_wire_1442[ 9 ] = fresh_wire_1439[ 9 ];
	assign fresh_wire_1442[ 10 ] = fresh_wire_1439[ 10 ];
	assign fresh_wire_1442[ 11 ] = fresh_wire_1439[ 11 ];
	assign fresh_wire_1442[ 12 ] = fresh_wire_1439[ 12 ];
	assign fresh_wire_1442[ 13 ] = fresh_wire_1439[ 13 ];
	assign fresh_wire_1442[ 14 ] = fresh_wire_1439[ 14 ];
	assign fresh_wire_1442[ 15 ] = fresh_wire_1439[ 15 ];
	assign fresh_wire_1444[ 0 ] = fresh_wire_1191[ 0 ];
	assign fresh_wire_1445[ 0 ] = fresh_wire_1374[ 0 ];
	assign fresh_wire_1445[ 1 ] = fresh_wire_1374[ 1 ];
	assign fresh_wire_1446[ 0 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1446[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1448[ 0 ] = fresh_wire_1301[ 0 ];
	assign fresh_wire_1449[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1449[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1450[ 0 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1450[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1452[ 0 ] = fresh_wire_1294[ 0 ];
	assign fresh_wire_1453[ 0 ] = fresh_wire_1447[ 0 ];
	assign fresh_wire_1453[ 1 ] = fresh_wire_1447[ 1 ];
	assign fresh_wire_1454[ 0 ] = fresh_wire_1451[ 0 ];
	assign fresh_wire_1454[ 1 ] = fresh_wire_1451[ 1 ];
	assign fresh_wire_1456[ 0 ] = fresh_wire_1289[ 0 ];
	assign fresh_wire_1457[ 0 ] = fresh_wire_1455[ 0 ];
	assign fresh_wire_1457[ 1 ] = fresh_wire_1455[ 1 ];
	assign fresh_wire_1458[ 0 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1458[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1460[ 0 ] = fresh_wire_1282[ 0 ];
	assign fresh_wire_1461[ 0 ] = fresh_wire_1459[ 0 ];
	assign fresh_wire_1461[ 1 ] = fresh_wire_1459[ 1 ];
	assign fresh_wire_1462[ 0 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1462[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1464[ 0 ] = fresh_wire_1270[ 0 ];
	assign fresh_wire_1465[ 0 ] = fresh_wire_1374[ 0 ];
	assign fresh_wire_1465[ 1 ] = fresh_wire_1374[ 1 ];
	assign fresh_wire_1466[ 0 ] = fresh_wire_1463[ 0 ];
	assign fresh_wire_1466[ 1 ] = fresh_wire_1463[ 1 ];
	assign fresh_wire_1468[ 0 ] = fresh_wire_1191[ 0 ];
	assign fresh_wire_1469[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1470[ 0 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1472[ 0 ] = fresh_wire_1289[ 0 ];
	assign fresh_wire_1473[ 0 ] = fresh_wire_1471[ 0 ];
	assign fresh_wire_1474[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1476[ 0 ] = fresh_wire_1282[ 0 ];
	assign fresh_wire_1477[ 0 ] = fresh_wire_1475[ 0 ];
	assign fresh_wire_1478[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1480[ 0 ] = fresh_wire_1270[ 0 ];
	assign fresh_wire_1481[ 0 ] = fresh_wire_1370[ 0 ];
	assign fresh_wire_1482[ 0 ] = fresh_wire_1479[ 0 ];
	assign fresh_wire_1484[ 0 ] = fresh_wire_1191[ 0 ];
	assign fresh_wire_1485[ 0 ] = fresh_wire_1366[ 0 ];
	assign fresh_wire_1486[ 0 ] = fresh_wire_1342[ 0 ];
	assign fresh_wire_1488[ 0 ] = fresh_wire_1301[ 0 ];
	assign fresh_wire_1489[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1490[ 0 ] = fresh_wire_1366[ 0 ];
	assign fresh_wire_1492[ 0 ] = fresh_wire_1294[ 0 ];
	assign fresh_wire_1493[ 0 ] = fresh_wire_1487[ 0 ];
	assign fresh_wire_1494[ 0 ] = fresh_wire_1491[ 0 ];
	assign fresh_wire_1496[ 0 ] = fresh_wire_1289[ 0 ];
	assign fresh_wire_1497[ 0 ] = fresh_wire_1495[ 0 ];
	assign fresh_wire_1498[ 0 ] = fresh_wire_1366[ 0 ];
	assign fresh_wire_1500[ 0 ] = fresh_wire_1282[ 0 ];
	assign fresh_wire_1501[ 0 ] = fresh_wire_1499[ 0 ];
	assign fresh_wire_1502[ 0 ] = fresh_wire_1342[ 0 ];
	assign fresh_wire_1504[ 0 ] = fresh_wire_1270[ 0 ];
	assign fresh_wire_1505[ 0 ] = fresh_wire_1366[ 0 ];
	assign fresh_wire_1506[ 0 ] = fresh_wire_1503[ 0 ];
	assign fresh_wire_1508[ 0 ] = fresh_wire_1191[ 0 ];
	assign fresh_wire_1509[ 0 ] = fresh_wire_1390[ 0 ];
	assign fresh_wire_1509[ 1 ] = fresh_wire_1390[ 1 ];
	assign fresh_wire_1509[ 2 ] = fresh_wire_1390[ 2 ];
	assign fresh_wire_1509[ 3 ] = fresh_wire_1390[ 3 ];
	assign fresh_wire_1509[ 4 ] = fresh_wire_1390[ 4 ];
	assign fresh_wire_1509[ 5 ] = fresh_wire_1390[ 5 ];
	assign fresh_wire_1509[ 6 ] = fresh_wire_1390[ 6 ];
	assign fresh_wire_1509[ 7 ] = fresh_wire_1390[ 7 ];
	assign fresh_wire_1509[ 8 ] = fresh_wire_1390[ 8 ];
	assign fresh_wire_1509[ 9 ] = fresh_wire_1390[ 9 ];
	assign fresh_wire_1509[ 10 ] = fresh_wire_1390[ 10 ];
	assign fresh_wire_1509[ 11 ] = fresh_wire_1390[ 11 ];
	assign fresh_wire_1509[ 12 ] = fresh_wire_1390[ 12 ];
	assign fresh_wire_1509[ 13 ] = fresh_wire_1390[ 13 ];
	assign fresh_wire_1509[ 14 ] = fresh_wire_1390[ 14 ];
	assign fresh_wire_1509[ 15 ] = fresh_wire_1390[ 15 ];
	assign fresh_wire_1510[ 0 ] = fresh_wire_1569[ 0 ];
	assign fresh_wire_1510[ 1 ] = fresh_wire_1569[ 1 ];
	assign fresh_wire_1510[ 2 ] = fresh_wire_1569[ 2 ];
	assign fresh_wire_1510[ 3 ] = fresh_wire_1569[ 3 ];
	assign fresh_wire_1510[ 4 ] = fresh_wire_1569[ 4 ];
	assign fresh_wire_1510[ 5 ] = fresh_wire_1569[ 5 ];
	assign fresh_wire_1510[ 6 ] = fresh_wire_1569[ 6 ];
	assign fresh_wire_1510[ 7 ] = fresh_wire_1569[ 7 ];
	assign fresh_wire_1510[ 8 ] = fresh_wire_1569[ 8 ];
	assign fresh_wire_1510[ 9 ] = fresh_wire_1569[ 9 ];
	assign fresh_wire_1510[ 10 ] = fresh_wire_1569[ 10 ];
	assign fresh_wire_1510[ 11 ] = fresh_wire_1569[ 11 ];
	assign fresh_wire_1510[ 12 ] = fresh_wire_1569[ 12 ];
	assign fresh_wire_1510[ 13 ] = fresh_wire_1569[ 13 ];
	assign fresh_wire_1510[ 14 ] = fresh_wire_1569[ 14 ];
	assign fresh_wire_1510[ 15 ] = fresh_wire_1569[ 15 ];
	assign fresh_wire_1512[ 0 ] = fresh_wire_1200[ 0 ];
	assign fresh_wire_1513[ 0 ] = fresh_wire_1390[ 0 ];
	assign fresh_wire_1513[ 1 ] = fresh_wire_1390[ 1 ];
	assign fresh_wire_1513[ 2 ] = fresh_wire_1390[ 2 ];
	assign fresh_wire_1513[ 3 ] = fresh_wire_1390[ 3 ];
	assign fresh_wire_1513[ 4 ] = fresh_wire_1390[ 4 ];
	assign fresh_wire_1513[ 5 ] = fresh_wire_1390[ 5 ];
	assign fresh_wire_1513[ 6 ] = fresh_wire_1390[ 6 ];
	assign fresh_wire_1513[ 7 ] = fresh_wire_1390[ 7 ];
	assign fresh_wire_1513[ 8 ] = fresh_wire_1390[ 8 ];
	assign fresh_wire_1513[ 9 ] = fresh_wire_1390[ 9 ];
	assign fresh_wire_1513[ 10 ] = fresh_wire_1390[ 10 ];
	assign fresh_wire_1513[ 11 ] = fresh_wire_1390[ 11 ];
	assign fresh_wire_1513[ 12 ] = fresh_wire_1390[ 12 ];
	assign fresh_wire_1513[ 13 ] = fresh_wire_1390[ 13 ];
	assign fresh_wire_1513[ 14 ] = fresh_wire_1390[ 14 ];
	assign fresh_wire_1513[ 15 ] = fresh_wire_1390[ 15 ];
	assign fresh_wire_1514[ 0 ] = fresh_wire_1153[ 0 ];
	assign fresh_wire_1514[ 1 ] = fresh_wire_1153[ 1 ];
	assign fresh_wire_1514[ 2 ] = fresh_wire_1153[ 2 ];
	assign fresh_wire_1514[ 3 ] = fresh_wire_1153[ 3 ];
	assign fresh_wire_1514[ 4 ] = fresh_wire_1153[ 4 ];
	assign fresh_wire_1514[ 5 ] = fresh_wire_1153[ 5 ];
	assign fresh_wire_1514[ 6 ] = fresh_wire_1153[ 6 ];
	assign fresh_wire_1514[ 7 ] = fresh_wire_1153[ 7 ];
	assign fresh_wire_1514[ 8 ] = fresh_wire_1153[ 8 ];
	assign fresh_wire_1514[ 9 ] = fresh_wire_1153[ 9 ];
	assign fresh_wire_1514[ 10 ] = fresh_wire_1153[ 10 ];
	assign fresh_wire_1514[ 11 ] = fresh_wire_1153[ 11 ];
	assign fresh_wire_1514[ 12 ] = fresh_wire_1153[ 12 ];
	assign fresh_wire_1514[ 13 ] = fresh_wire_1153[ 13 ];
	assign fresh_wire_1514[ 14 ] = fresh_wire_1153[ 14 ];
	assign fresh_wire_1514[ 15 ] = fresh_wire_1153[ 15 ];
	assign fresh_wire_1516[ 0 ] = fresh_wire_1206[ 0 ];
	assign fresh_wire_1517[ 0 ] = fresh_wire_1511[ 0 ];
	assign fresh_wire_1517[ 1 ] = fresh_wire_1511[ 1 ];
	assign fresh_wire_1517[ 2 ] = fresh_wire_1511[ 2 ];
	assign fresh_wire_1517[ 3 ] = fresh_wire_1511[ 3 ];
	assign fresh_wire_1517[ 4 ] = fresh_wire_1511[ 4 ];
	assign fresh_wire_1517[ 5 ] = fresh_wire_1511[ 5 ];
	assign fresh_wire_1517[ 6 ] = fresh_wire_1511[ 6 ];
	assign fresh_wire_1517[ 7 ] = fresh_wire_1511[ 7 ];
	assign fresh_wire_1517[ 8 ] = fresh_wire_1511[ 8 ];
	assign fresh_wire_1517[ 9 ] = fresh_wire_1511[ 9 ];
	assign fresh_wire_1517[ 10 ] = fresh_wire_1511[ 10 ];
	assign fresh_wire_1517[ 11 ] = fresh_wire_1511[ 11 ];
	assign fresh_wire_1517[ 12 ] = fresh_wire_1511[ 12 ];
	assign fresh_wire_1517[ 13 ] = fresh_wire_1511[ 13 ];
	assign fresh_wire_1517[ 14 ] = fresh_wire_1511[ 14 ];
	assign fresh_wire_1517[ 15 ] = fresh_wire_1511[ 15 ];
	assign fresh_wire_1518[ 0 ] = fresh_wire_1515[ 0 ];
	assign fresh_wire_1518[ 1 ] = fresh_wire_1515[ 1 ];
	assign fresh_wire_1518[ 2 ] = fresh_wire_1515[ 2 ];
	assign fresh_wire_1518[ 3 ] = fresh_wire_1515[ 3 ];
	assign fresh_wire_1518[ 4 ] = fresh_wire_1515[ 4 ];
	assign fresh_wire_1518[ 5 ] = fresh_wire_1515[ 5 ];
	assign fresh_wire_1518[ 6 ] = fresh_wire_1515[ 6 ];
	assign fresh_wire_1518[ 7 ] = fresh_wire_1515[ 7 ];
	assign fresh_wire_1518[ 8 ] = fresh_wire_1515[ 8 ];
	assign fresh_wire_1518[ 9 ] = fresh_wire_1515[ 9 ];
	assign fresh_wire_1518[ 10 ] = fresh_wire_1515[ 10 ];
	assign fresh_wire_1518[ 11 ] = fresh_wire_1515[ 11 ];
	assign fresh_wire_1518[ 12 ] = fresh_wire_1515[ 12 ];
	assign fresh_wire_1518[ 13 ] = fresh_wire_1515[ 13 ];
	assign fresh_wire_1518[ 14 ] = fresh_wire_1515[ 14 ];
	assign fresh_wire_1518[ 15 ] = fresh_wire_1515[ 15 ];
	assign fresh_wire_1520[ 0 ] = fresh_wire_1203[ 0 ];
	assign fresh_wire_1521[ 0 ] = fresh_wire_1148[ 0 ];
	assign fresh_wire_1521[ 1 ] = fresh_wire_1148[ 1 ];
	assign fresh_wire_1521[ 2 ] = fresh_wire_1148[ 2 ];
	assign fresh_wire_1521[ 3 ] = fresh_wire_1148[ 3 ];
	assign fresh_wire_1521[ 4 ] = fresh_wire_1148[ 4 ];
	assign fresh_wire_1521[ 5 ] = fresh_wire_1148[ 5 ];
	assign fresh_wire_1521[ 6 ] = fresh_wire_1148[ 6 ];
	assign fresh_wire_1521[ 7 ] = fresh_wire_1148[ 7 ];
	assign fresh_wire_1521[ 8 ] = fresh_wire_1148[ 8 ];
	assign fresh_wire_1521[ 9 ] = fresh_wire_1148[ 9 ];
	assign fresh_wire_1521[ 10 ] = fresh_wire_1148[ 10 ];
	assign fresh_wire_1521[ 11 ] = fresh_wire_1148[ 11 ];
	assign fresh_wire_1521[ 12 ] = fresh_wire_1148[ 12 ];
	assign fresh_wire_1521[ 13 ] = fresh_wire_1148[ 13 ];
	assign fresh_wire_1521[ 14 ] = fresh_wire_1148[ 14 ];
	assign fresh_wire_1521[ 15 ] = fresh_wire_1148[ 15 ];
	assign fresh_wire_1522[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1522[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1522[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1522[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1522[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1522[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1522[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1522[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1522[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1522[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1522[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1522[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1522[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1522[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1522[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1522[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1524[ 0 ] = fresh_wire_1233[ 0 ];
	assign fresh_wire_1525[ 0 ] = fresh_wire_1386[ 0 ];
	assign fresh_wire_1525[ 1 ] = fresh_wire_1386[ 1 ];
	assign fresh_wire_1525[ 2 ] = fresh_wire_1386[ 2 ];
	assign fresh_wire_1525[ 3 ] = fresh_wire_1386[ 3 ];
	assign fresh_wire_1525[ 4 ] = fresh_wire_1386[ 4 ];
	assign fresh_wire_1525[ 5 ] = fresh_wire_1386[ 5 ];
	assign fresh_wire_1525[ 6 ] = fresh_wire_1386[ 6 ];
	assign fresh_wire_1525[ 7 ] = fresh_wire_1386[ 7 ];
	assign fresh_wire_1525[ 8 ] = fresh_wire_1386[ 8 ];
	assign fresh_wire_1525[ 9 ] = fresh_wire_1386[ 9 ];
	assign fresh_wire_1525[ 10 ] = fresh_wire_1386[ 10 ];
	assign fresh_wire_1525[ 11 ] = fresh_wire_1386[ 11 ];
	assign fresh_wire_1525[ 12 ] = fresh_wire_1386[ 12 ];
	assign fresh_wire_1525[ 13 ] = fresh_wire_1386[ 13 ];
	assign fresh_wire_1525[ 14 ] = fresh_wire_1386[ 14 ];
	assign fresh_wire_1525[ 15 ] = fresh_wire_1386[ 15 ];
	assign fresh_wire_1526[ 0 ] = fresh_wire_1523[ 0 ];
	assign fresh_wire_1526[ 1 ] = fresh_wire_1523[ 1 ];
	assign fresh_wire_1526[ 2 ] = fresh_wire_1523[ 2 ];
	assign fresh_wire_1526[ 3 ] = fresh_wire_1523[ 3 ];
	assign fresh_wire_1526[ 4 ] = fresh_wire_1523[ 4 ];
	assign fresh_wire_1526[ 5 ] = fresh_wire_1523[ 5 ];
	assign fresh_wire_1526[ 6 ] = fresh_wire_1523[ 6 ];
	assign fresh_wire_1526[ 7 ] = fresh_wire_1523[ 7 ];
	assign fresh_wire_1526[ 8 ] = fresh_wire_1523[ 8 ];
	assign fresh_wire_1526[ 9 ] = fresh_wire_1523[ 9 ];
	assign fresh_wire_1526[ 10 ] = fresh_wire_1523[ 10 ];
	assign fresh_wire_1526[ 11 ] = fresh_wire_1523[ 11 ];
	assign fresh_wire_1526[ 12 ] = fresh_wire_1523[ 12 ];
	assign fresh_wire_1526[ 13 ] = fresh_wire_1523[ 13 ];
	assign fresh_wire_1526[ 14 ] = fresh_wire_1523[ 14 ];
	assign fresh_wire_1526[ 15 ] = fresh_wire_1523[ 15 ];
	assign fresh_wire_1528[ 0 ] = fresh_wire_1206[ 0 ];
	assign fresh_wire_1529[ 0 ] = fresh_wire_1386[ 0 ];
	assign fresh_wire_1529[ 1 ] = fresh_wire_1386[ 1 ];
	assign fresh_wire_1529[ 2 ] = fresh_wire_1386[ 2 ];
	assign fresh_wire_1529[ 3 ] = fresh_wire_1386[ 3 ];
	assign fresh_wire_1529[ 4 ] = fresh_wire_1386[ 4 ];
	assign fresh_wire_1529[ 5 ] = fresh_wire_1386[ 5 ];
	assign fresh_wire_1529[ 6 ] = fresh_wire_1386[ 6 ];
	assign fresh_wire_1529[ 7 ] = fresh_wire_1386[ 7 ];
	assign fresh_wire_1529[ 8 ] = fresh_wire_1386[ 8 ];
	assign fresh_wire_1529[ 9 ] = fresh_wire_1386[ 9 ];
	assign fresh_wire_1529[ 10 ] = fresh_wire_1386[ 10 ];
	assign fresh_wire_1529[ 11 ] = fresh_wire_1386[ 11 ];
	assign fresh_wire_1529[ 12 ] = fresh_wire_1386[ 12 ];
	assign fresh_wire_1529[ 13 ] = fresh_wire_1386[ 13 ];
	assign fresh_wire_1529[ 14 ] = fresh_wire_1386[ 14 ];
	assign fresh_wire_1529[ 15 ] = fresh_wire_1386[ 15 ];
	assign fresh_wire_1530[ 0 ] = fresh_wire_1527[ 0 ];
	assign fresh_wire_1530[ 1 ] = fresh_wire_1527[ 1 ];
	assign fresh_wire_1530[ 2 ] = fresh_wire_1527[ 2 ];
	assign fresh_wire_1530[ 3 ] = fresh_wire_1527[ 3 ];
	assign fresh_wire_1530[ 4 ] = fresh_wire_1527[ 4 ];
	assign fresh_wire_1530[ 5 ] = fresh_wire_1527[ 5 ];
	assign fresh_wire_1530[ 6 ] = fresh_wire_1527[ 6 ];
	assign fresh_wire_1530[ 7 ] = fresh_wire_1527[ 7 ];
	assign fresh_wire_1530[ 8 ] = fresh_wire_1527[ 8 ];
	assign fresh_wire_1530[ 9 ] = fresh_wire_1527[ 9 ];
	assign fresh_wire_1530[ 10 ] = fresh_wire_1527[ 10 ];
	assign fresh_wire_1530[ 11 ] = fresh_wire_1527[ 11 ];
	assign fresh_wire_1530[ 12 ] = fresh_wire_1527[ 12 ];
	assign fresh_wire_1530[ 13 ] = fresh_wire_1527[ 13 ];
	assign fresh_wire_1530[ 14 ] = fresh_wire_1527[ 14 ];
	assign fresh_wire_1530[ 15 ] = fresh_wire_1527[ 15 ];
	assign fresh_wire_1532[ 0 ] = fresh_wire_1203[ 0 ];
	assign fresh_wire_1533[ 0 ] = fresh_wire_1158[ 0 ];
	assign fresh_wire_1533[ 1 ] = fresh_wire_1158[ 1 ];
	assign fresh_wire_1533[ 2 ] = fresh_wire_1158[ 2 ];
	assign fresh_wire_1533[ 3 ] = fresh_wire_1158[ 3 ];
	assign fresh_wire_1533[ 4 ] = fresh_wire_1158[ 4 ];
	assign fresh_wire_1533[ 5 ] = fresh_wire_1158[ 5 ];
	assign fresh_wire_1533[ 6 ] = fresh_wire_1158[ 6 ];
	assign fresh_wire_1533[ 7 ] = fresh_wire_1158[ 7 ];
	assign fresh_wire_1533[ 8 ] = fresh_wire_1158[ 8 ];
	assign fresh_wire_1533[ 9 ] = fresh_wire_1158[ 9 ];
	assign fresh_wire_1533[ 10 ] = fresh_wire_1158[ 10 ];
	assign fresh_wire_1533[ 11 ] = fresh_wire_1158[ 11 ];
	assign fresh_wire_1533[ 12 ] = fresh_wire_1158[ 12 ];
	assign fresh_wire_1533[ 13 ] = fresh_wire_1158[ 13 ];
	assign fresh_wire_1533[ 14 ] = fresh_wire_1158[ 14 ];
	assign fresh_wire_1533[ 15 ] = fresh_wire_1158[ 15 ];
	assign fresh_wire_1534[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1534[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1534[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1534[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1534[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1534[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1534[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1534[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1534[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1534[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1534[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1534[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1534[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1534[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1534[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1534[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1536[ 0 ] = fresh_wire_1236[ 0 ];
	assign fresh_wire_1537[ 0 ] = fresh_wire_1382[ 0 ];
	assign fresh_wire_1537[ 1 ] = fresh_wire_1382[ 1 ];
	assign fresh_wire_1537[ 2 ] = fresh_wire_1382[ 2 ];
	assign fresh_wire_1537[ 3 ] = fresh_wire_1382[ 3 ];
	assign fresh_wire_1537[ 4 ] = fresh_wire_1382[ 4 ];
	assign fresh_wire_1537[ 5 ] = fresh_wire_1382[ 5 ];
	assign fresh_wire_1537[ 6 ] = fresh_wire_1382[ 6 ];
	assign fresh_wire_1537[ 7 ] = fresh_wire_1382[ 7 ];
	assign fresh_wire_1537[ 8 ] = fresh_wire_1382[ 8 ];
	assign fresh_wire_1537[ 9 ] = fresh_wire_1382[ 9 ];
	assign fresh_wire_1537[ 10 ] = fresh_wire_1382[ 10 ];
	assign fresh_wire_1537[ 11 ] = fresh_wire_1382[ 11 ];
	assign fresh_wire_1537[ 12 ] = fresh_wire_1382[ 12 ];
	assign fresh_wire_1537[ 13 ] = fresh_wire_1382[ 13 ];
	assign fresh_wire_1537[ 14 ] = fresh_wire_1382[ 14 ];
	assign fresh_wire_1537[ 15 ] = fresh_wire_1382[ 15 ];
	assign fresh_wire_1538[ 0 ] = fresh_wire_1535[ 0 ];
	assign fresh_wire_1538[ 1 ] = fresh_wire_1535[ 1 ];
	assign fresh_wire_1538[ 2 ] = fresh_wire_1535[ 2 ];
	assign fresh_wire_1538[ 3 ] = fresh_wire_1535[ 3 ];
	assign fresh_wire_1538[ 4 ] = fresh_wire_1535[ 4 ];
	assign fresh_wire_1538[ 5 ] = fresh_wire_1535[ 5 ];
	assign fresh_wire_1538[ 6 ] = fresh_wire_1535[ 6 ];
	assign fresh_wire_1538[ 7 ] = fresh_wire_1535[ 7 ];
	assign fresh_wire_1538[ 8 ] = fresh_wire_1535[ 8 ];
	assign fresh_wire_1538[ 9 ] = fresh_wire_1535[ 9 ];
	assign fresh_wire_1538[ 10 ] = fresh_wire_1535[ 10 ];
	assign fresh_wire_1538[ 11 ] = fresh_wire_1535[ 11 ];
	assign fresh_wire_1538[ 12 ] = fresh_wire_1535[ 12 ];
	assign fresh_wire_1538[ 13 ] = fresh_wire_1535[ 13 ];
	assign fresh_wire_1538[ 14 ] = fresh_wire_1535[ 14 ];
	assign fresh_wire_1538[ 15 ] = fresh_wire_1535[ 15 ];
	assign fresh_wire_1540[ 0 ] = fresh_wire_1200[ 0 ];
	assign fresh_wire_1541[ 0 ] = fresh_wire_1539[ 0 ];
	assign fresh_wire_1541[ 1 ] = fresh_wire_1539[ 1 ];
	assign fresh_wire_1541[ 2 ] = fresh_wire_1539[ 2 ];
	assign fresh_wire_1541[ 3 ] = fresh_wire_1539[ 3 ];
	assign fresh_wire_1541[ 4 ] = fresh_wire_1539[ 4 ];
	assign fresh_wire_1541[ 5 ] = fresh_wire_1539[ 5 ];
	assign fresh_wire_1541[ 6 ] = fresh_wire_1539[ 6 ];
	assign fresh_wire_1541[ 7 ] = fresh_wire_1539[ 7 ];
	assign fresh_wire_1541[ 8 ] = fresh_wire_1539[ 8 ];
	assign fresh_wire_1541[ 9 ] = fresh_wire_1539[ 9 ];
	assign fresh_wire_1541[ 10 ] = fresh_wire_1539[ 10 ];
	assign fresh_wire_1541[ 11 ] = fresh_wire_1539[ 11 ];
	assign fresh_wire_1541[ 12 ] = fresh_wire_1539[ 12 ];
	assign fresh_wire_1541[ 13 ] = fresh_wire_1539[ 13 ];
	assign fresh_wire_1541[ 14 ] = fresh_wire_1539[ 14 ];
	assign fresh_wire_1541[ 15 ] = fresh_wire_1539[ 15 ];
	assign fresh_wire_1542[ 0 ] = fresh_wire_1382[ 0 ];
	assign fresh_wire_1542[ 1 ] = fresh_wire_1382[ 1 ];
	assign fresh_wire_1542[ 2 ] = fresh_wire_1382[ 2 ];
	assign fresh_wire_1542[ 3 ] = fresh_wire_1382[ 3 ];
	assign fresh_wire_1542[ 4 ] = fresh_wire_1382[ 4 ];
	assign fresh_wire_1542[ 5 ] = fresh_wire_1382[ 5 ];
	assign fresh_wire_1542[ 6 ] = fresh_wire_1382[ 6 ];
	assign fresh_wire_1542[ 7 ] = fresh_wire_1382[ 7 ];
	assign fresh_wire_1542[ 8 ] = fresh_wire_1382[ 8 ];
	assign fresh_wire_1542[ 9 ] = fresh_wire_1382[ 9 ];
	assign fresh_wire_1542[ 10 ] = fresh_wire_1382[ 10 ];
	assign fresh_wire_1542[ 11 ] = fresh_wire_1382[ 11 ];
	assign fresh_wire_1542[ 12 ] = fresh_wire_1382[ 12 ];
	assign fresh_wire_1542[ 13 ] = fresh_wire_1382[ 13 ];
	assign fresh_wire_1542[ 14 ] = fresh_wire_1382[ 14 ];
	assign fresh_wire_1542[ 15 ] = fresh_wire_1382[ 15 ];
	assign fresh_wire_1544[ 0 ] = fresh_wire_1203[ 0 ];
	assign fresh_wire_1545[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1546[ 0 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1548[ 0 ] = fresh_wire_1194[ 0 ];
	assign fresh_wire_1549[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1550[ 0 ] = fresh_wire_1547[ 0 ];
	assign fresh_wire_1552[ 0 ] = fresh_wire_1191[ 0 ];
	assign fresh_wire_1553[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1554[ 0 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1556[ 0 ] = fresh_wire_1197[ 0 ];
	assign fresh_wire_1557[ 0 ] = fresh_wire_1555[ 0 ];
	assign fresh_wire_1558[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1560[ 0 ] = fresh_wire_1194[ 0 ];
	assign fresh_wire_1561[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1562[ 0 ] = fresh_wire_1559[ 0 ];
	assign fresh_wire_1564[ 0 ] = fresh_wire_1191[ 0 ];
	assign fresh_wire_1565[ 0 ] = fresh_wire_1390[ 0 ];
	assign fresh_wire_1565[ 1 ] = fresh_wire_1390[ 1 ];
	assign fresh_wire_1565[ 2 ] = fresh_wire_1390[ 2 ];
	assign fresh_wire_1565[ 3 ] = fresh_wire_1390[ 3 ];
	assign fresh_wire_1565[ 4 ] = fresh_wire_1390[ 4 ];
	assign fresh_wire_1565[ 5 ] = fresh_wire_1390[ 5 ];
	assign fresh_wire_1565[ 6 ] = fresh_wire_1390[ 6 ];
	assign fresh_wire_1565[ 7 ] = fresh_wire_1390[ 7 ];
	assign fresh_wire_1565[ 8 ] = fresh_wire_1390[ 8 ];
	assign fresh_wire_1565[ 9 ] = fresh_wire_1390[ 9 ];
	assign fresh_wire_1565[ 10 ] = fresh_wire_1390[ 10 ];
	assign fresh_wire_1565[ 11 ] = fresh_wire_1390[ 11 ];
	assign fresh_wire_1565[ 12 ] = fresh_wire_1390[ 12 ];
	assign fresh_wire_1565[ 13 ] = fresh_wire_1390[ 13 ];
	assign fresh_wire_1565[ 14 ] = fresh_wire_1390[ 14 ];
	assign fresh_wire_1565[ 15 ] = fresh_wire_1390[ 15 ];
	assign fresh_wire_1567[ 0 ] = fresh_wire_1566[ 0 ];
	assign fresh_wire_1567[ 1 ] = fresh_wire_1566[ 1 ];
	assign fresh_wire_1567[ 2 ] = fresh_wire_1566[ 2 ];
	assign fresh_wire_1567[ 3 ] = fresh_wire_1566[ 3 ];
	assign fresh_wire_1567[ 4 ] = fresh_wire_1566[ 4 ];
	assign fresh_wire_1567[ 5 ] = fresh_wire_1566[ 5 ];
	assign fresh_wire_1567[ 6 ] = fresh_wire_1566[ 6 ];
	assign fresh_wire_1567[ 7 ] = fresh_wire_1566[ 7 ];
	assign fresh_wire_1567[ 8 ] = fresh_wire_1566[ 8 ];
	assign fresh_wire_1567[ 9 ] = fresh_wire_1566[ 9 ];
	assign fresh_wire_1567[ 10 ] = fresh_wire_1566[ 10 ];
	assign fresh_wire_1567[ 11 ] = fresh_wire_1566[ 11 ];
	assign fresh_wire_1567[ 12 ] = fresh_wire_1566[ 12 ];
	assign fresh_wire_1567[ 13 ] = fresh_wire_1566[ 13 ];
	assign fresh_wire_1567[ 14 ] = fresh_wire_1566[ 14 ];
	assign fresh_wire_1567[ 15 ] = fresh_wire_1566[ 15 ];
	assign fresh_wire_1567[ 16 ] = fresh_wire_1566[ 16 ];
	assign fresh_wire_1567[ 17 ] = fresh_wire_1566[ 17 ];
	assign fresh_wire_1567[ 18 ] = fresh_wire_1566[ 18 ];
	assign fresh_wire_1567[ 19 ] = fresh_wire_1566[ 19 ];
	assign fresh_wire_1567[ 20 ] = fresh_wire_1566[ 20 ];
	assign fresh_wire_1567[ 21 ] = fresh_wire_1566[ 21 ];
	assign fresh_wire_1567[ 22 ] = fresh_wire_1566[ 22 ];
	assign fresh_wire_1567[ 23 ] = fresh_wire_1566[ 23 ];
	assign fresh_wire_1567[ 24 ] = fresh_wire_1566[ 24 ];
	assign fresh_wire_1567[ 25 ] = fresh_wire_1566[ 25 ];
	assign fresh_wire_1567[ 26 ] = fresh_wire_1566[ 26 ];
	assign fresh_wire_1567[ 27 ] = fresh_wire_1566[ 27 ];
	assign fresh_wire_1567[ 28 ] = fresh_wire_1566[ 28 ];
	assign fresh_wire_1567[ 29 ] = fresh_wire_1566[ 29 ];
	assign fresh_wire_1567[ 30 ] = fresh_wire_1566[ 30 ];
	assign fresh_wire_1567[ 31 ] = fresh_wire_1566[ 31 ];
	assign fresh_wire_1568[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 1 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1568[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 16 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 17 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 18 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 19 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 20 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 21 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 22 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 23 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 24 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 25 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 26 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 27 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 28 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 29 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 30 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1568[ 31 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1570[ 0 ] = fresh_wire_1911[ 0 ];
	assign fresh_wire_1570[ 1 ] = fresh_wire_1911[ 1 ];
	assign fresh_wire_1570[ 2 ] = fresh_wire_1911[ 2 ];
	assign fresh_wire_1570[ 3 ] = fresh_wire_1911[ 3 ];
	assign fresh_wire_1570[ 4 ] = fresh_wire_1911[ 4 ];
	assign fresh_wire_1570[ 5 ] = fresh_wire_1911[ 5 ];
	assign fresh_wire_1570[ 6 ] = fresh_wire_1911[ 6 ];
	assign fresh_wire_1570[ 7 ] = fresh_wire_1911[ 7 ];
	assign fresh_wire_1570[ 8 ] = fresh_wire_1911[ 8 ];
	assign fresh_wire_1570[ 9 ] = fresh_wire_1911[ 9 ];
	assign fresh_wire_1570[ 10 ] = fresh_wire_1911[ 10 ];
	assign fresh_wire_1570[ 11 ] = fresh_wire_1911[ 11 ];
	assign fresh_wire_1570[ 12 ] = fresh_wire_1911[ 12 ];
	assign fresh_wire_1570[ 13 ] = fresh_wire_1911[ 13 ];
	assign fresh_wire_1570[ 14 ] = fresh_wire_1911[ 14 ];
	assign fresh_wire_1570[ 15 ] = fresh_wire_1911[ 15 ];
	assign fresh_wire_1570[ 16 ] = fresh_wire_2009[ 0 ];
	assign fresh_wire_1570[ 17 ] = fresh_wire_2009[ 1 ];
	assign fresh_wire_1570[ 18 ] = fresh_wire_2009[ 2 ];
	assign fresh_wire_1570[ 19 ] = fresh_wire_2009[ 3 ];
	assign fresh_wire_1570[ 20 ] = fresh_wire_2009[ 4 ];
	assign fresh_wire_1570[ 21 ] = fresh_wire_2009[ 5 ];
	assign fresh_wire_1570[ 22 ] = fresh_wire_2009[ 6 ];
	assign fresh_wire_1570[ 23 ] = fresh_wire_2009[ 7 ];
	assign fresh_wire_1570[ 24 ] = fresh_wire_2009[ 8 ];
	assign fresh_wire_1570[ 25 ] = fresh_wire_2009[ 9 ];
	assign fresh_wire_1570[ 26 ] = fresh_wire_2009[ 10 ];
	assign fresh_wire_1570[ 27 ] = fresh_wire_2009[ 11 ];
	assign fresh_wire_1570[ 28 ] = fresh_wire_2009[ 12 ];
	assign fresh_wire_1570[ 29 ] = fresh_wire_2009[ 13 ];
	assign fresh_wire_1570[ 30 ] = fresh_wire_2009[ 14 ];
	assign fresh_wire_1570[ 31 ] = fresh_wire_2009[ 15 ];
	assign fresh_wire_1571[ 0 ] = fresh_wire_1686[ 0 ];
	assign fresh_wire_1571[ 1 ] = fresh_wire_1686[ 1 ];
	assign fresh_wire_1571[ 2 ] = fresh_wire_1686[ 2 ];
	assign fresh_wire_1571[ 3 ] = fresh_wire_1686[ 3 ];
	assign fresh_wire_1571[ 4 ] = fresh_wire_1686[ 4 ];
	assign fresh_wire_1571[ 5 ] = fresh_wire_1686[ 5 ];
	assign fresh_wire_1571[ 6 ] = fresh_wire_1686[ 6 ];
	assign fresh_wire_1571[ 7 ] = fresh_wire_1686[ 7 ];
	assign fresh_wire_1571[ 8 ] = fresh_wire_1686[ 8 ];
	assign fresh_wire_1571[ 9 ] = fresh_wire_1686[ 9 ];
	assign fresh_wire_1571[ 10 ] = fresh_wire_1686[ 10 ];
	assign fresh_wire_1571[ 11 ] = fresh_wire_1686[ 11 ];
	assign fresh_wire_1571[ 12 ] = fresh_wire_1686[ 12 ];
	assign fresh_wire_1571[ 13 ] = fresh_wire_1686[ 13 ];
	assign fresh_wire_1571[ 14 ] = fresh_wire_1686[ 14 ];
	assign fresh_wire_1571[ 15 ] = fresh_wire_1686[ 15 ];
	assign fresh_wire_1571[ 16 ] = fresh_wire_1686[ 16 ];
	assign fresh_wire_1571[ 17 ] = fresh_wire_1686[ 17 ];
	assign fresh_wire_1571[ 18 ] = fresh_wire_1686[ 18 ];
	assign fresh_wire_1571[ 19 ] = fresh_wire_1686[ 19 ];
	assign fresh_wire_1571[ 20 ] = fresh_wire_1686[ 20 ];
	assign fresh_wire_1571[ 21 ] = fresh_wire_1686[ 21 ];
	assign fresh_wire_1571[ 22 ] = fresh_wire_1686[ 22 ];
	assign fresh_wire_1571[ 23 ] = fresh_wire_1686[ 23 ];
	assign fresh_wire_1571[ 24 ] = fresh_wire_1686[ 24 ];
	assign fresh_wire_1571[ 25 ] = fresh_wire_1686[ 25 ];
	assign fresh_wire_1571[ 26 ] = fresh_wire_1686[ 26 ];
	assign fresh_wire_1571[ 27 ] = fresh_wire_1686[ 27 ];
	assign fresh_wire_1571[ 28 ] = fresh_wire_1686[ 28 ];
	assign fresh_wire_1571[ 29 ] = fresh_wire_1686[ 29 ];
	assign fresh_wire_1571[ 30 ] = fresh_wire_1686[ 30 ];
	assign fresh_wire_1571[ 31 ] = fresh_wire_1686[ 31 ];
	assign fresh_wire_1573[ 0 ] = fresh_wire_1188[ 0 ];
	assign fresh_wire_1574[ 0 ] = fresh_wire_1164[ 0 ];
	assign fresh_wire_1574[ 1 ] = fresh_wire_1164[ 1 ];
	assign fresh_wire_1574[ 2 ] = fresh_wire_1164[ 2 ];
	assign fresh_wire_1574[ 3 ] = fresh_wire_1164[ 3 ];
	assign fresh_wire_1574[ 4 ] = fresh_wire_1164[ 4 ];
	assign fresh_wire_1574[ 5 ] = fresh_wire_1164[ 5 ];
	assign fresh_wire_1574[ 6 ] = fresh_wire_1164[ 6 ];
	assign fresh_wire_1574[ 7 ] = fresh_wire_1164[ 7 ];
	assign fresh_wire_1574[ 8 ] = fresh_wire_1164[ 8 ];
	assign fresh_wire_1574[ 9 ] = fresh_wire_1164[ 9 ];
	assign fresh_wire_1574[ 10 ] = fresh_wire_1164[ 10 ];
	assign fresh_wire_1574[ 11 ] = fresh_wire_1164[ 11 ];
	assign fresh_wire_1574[ 12 ] = fresh_wire_1164[ 12 ];
	assign fresh_wire_1574[ 13 ] = fresh_wire_1164[ 13 ];
	assign fresh_wire_1574[ 14 ] = fresh_wire_1164[ 14 ];
	assign fresh_wire_1574[ 15 ] = fresh_wire_1164[ 15 ];
	assign fresh_wire_1575[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1575[ 1 ] = fresh_wire_1578[ 0 ];
	assign fresh_wire_1575[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1575[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1575[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1575[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1575[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1575[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1575[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1575[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1575[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1575[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1575[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1575[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1575[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1575[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1577[ 0 ] = fresh_wire_1215[ 0 ];
	assign fresh_wire_1579[ 0 ] = fresh_wire_1850[ 0 ];
	assign fresh_wire_1579[ 1 ] = fresh_wire_1850[ 1 ];
	assign fresh_wire_1579[ 2 ] = fresh_wire_1850[ 2 ];
	assign fresh_wire_1579[ 3 ] = fresh_wire_1850[ 3 ];
	assign fresh_wire_1579[ 4 ] = fresh_wire_1850[ 4 ];
	assign fresh_wire_1579[ 5 ] = fresh_wire_1850[ 5 ];
	assign fresh_wire_1579[ 6 ] = fresh_wire_1850[ 6 ];
	assign fresh_wire_1579[ 7 ] = fresh_wire_1850[ 7 ];
	assign fresh_wire_1579[ 8 ] = fresh_wire_1850[ 8 ];
	assign fresh_wire_1579[ 9 ] = fresh_wire_1850[ 9 ];
	assign fresh_wire_1579[ 10 ] = fresh_wire_1850[ 10 ];
	assign fresh_wire_1579[ 11 ] = fresh_wire_1850[ 11 ];
	assign fresh_wire_1579[ 12 ] = fresh_wire_1850[ 12 ];
	assign fresh_wire_1579[ 13 ] = fresh_wire_1850[ 13 ];
	assign fresh_wire_1579[ 14 ] = fresh_wire_1850[ 14 ];
	assign fresh_wire_1579[ 15 ] = fresh_wire_1850[ 15 ];
	assign fresh_wire_1580[ 0 ] = fresh_wire_1351[ 0 ];
	assign fresh_wire_1580[ 1 ] = fresh_wire_1351[ 1 ];
	assign fresh_wire_1580[ 2 ] = fresh_wire_1351[ 2 ];
	assign fresh_wire_1580[ 3 ] = fresh_wire_1351[ 3 ];
	assign fresh_wire_1580[ 4 ] = fresh_wire_1351[ 4 ];
	assign fresh_wire_1580[ 5 ] = fresh_wire_1351[ 5 ];
	assign fresh_wire_1580[ 6 ] = fresh_wire_1351[ 6 ];
	assign fresh_wire_1580[ 7 ] = fresh_wire_1351[ 7 ];
	assign fresh_wire_1580[ 8 ] = fresh_wire_1351[ 8 ];
	assign fresh_wire_1580[ 9 ] = fresh_wire_1351[ 9 ];
	assign fresh_wire_1580[ 10 ] = fresh_wire_1351[ 10 ];
	assign fresh_wire_1580[ 11 ] = fresh_wire_1351[ 11 ];
	assign fresh_wire_1580[ 12 ] = fresh_wire_1351[ 12 ];
	assign fresh_wire_1580[ 13 ] = fresh_wire_1351[ 13 ];
	assign fresh_wire_1580[ 14 ] = fresh_wire_1351[ 14 ];
	assign fresh_wire_1580[ 15 ] = fresh_wire_1351[ 15 ];
	assign fresh_wire_1582[ 0 ] = fresh_wire_1230[ 0 ];
	assign fresh_wire_1583[ 0 ] = fresh_wire_1638[ 0 ];
	assign fresh_wire_1583[ 1 ] = fresh_wire_1638[ 1 ];
	assign fresh_wire_1584[ 0 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1584[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1586[ 0 ] = fresh_wire_1398[ 0 ];
	assign fresh_wire_1587[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1589[ 0 ] = fresh_wire_1394[ 0 ];
	assign fresh_wire_1590[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1592[ 0 ] = fresh_wire_1398[ 0 ];
	assign fresh_wire_1593[ 0 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1595[ 0 ] = fresh_wire_1638[ 0 ];
	assign fresh_wire_1595[ 1 ] = fresh_wire_1638[ 1 ];
	assign fresh_wire_1596[ 0 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1596[ 1 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1598[ 0 ] = fresh_wire_1638[ 0 ];
	assign fresh_wire_1598[ 1 ] = fresh_wire_1638[ 1 ];
	assign fresh_wire_1599[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1599[ 1 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1601[ 0 ] = fresh_wire_1394[ 0 ];
	assign fresh_wire_1602[ 0 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1604[ 0 ] = fresh_wire_1638[ 0 ];
	assign fresh_wire_1604[ 1 ] = fresh_wire_1638[ 1 ];
	assign fresh_wire_1605[ 0 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1605[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1607[ 0 ] = fresh_wire_1638[ 0 ];
	assign fresh_wire_1607[ 1 ] = fresh_wire_1638[ 1 ];
	assign fresh_wire_1608[ 0 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1608[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1610[ 0 ] = fresh_wire_1588[ 0 ];
	assign fresh_wire_1612[ 0 ] = fresh_wire_1611[ 0 ];
	assign fresh_wire_1613[ 0 ] = fresh_wire_1616[ 0 ];
	assign fresh_wire_1615[ 0 ] = fresh_wire_1591[ 0 ];
	assign fresh_wire_1617[ 0 ] = fresh_wire_2290[ 0 ];
	assign fresh_wire_1618[ 0 ] = fresh_wire_1621[ 0 ];
	assign fresh_wire_1620[ 0 ] = fresh_wire_1614[ 0 ];
	assign fresh_wire_1622[ 0 ] = fresh_wire_2291[ 0 ];
	assign fresh_wire_1623[ 0 ] = fresh_wire_1626[ 0 ];
	assign fresh_wire_1625[ 0 ] = fresh_wire_1594[ 0 ];
	assign fresh_wire_1627[ 0 ] = fresh_wire_2292[ 0 ];
	assign fresh_wire_1628[ 0 ] = fresh_wire_1631[ 0 ];
	assign fresh_wire_1630[ 0 ] = fresh_wire_1588[ 0 ];
	assign fresh_wire_1632[ 0 ] = fresh_wire_2293[ 0 ];
	assign fresh_wire_1633[ 0 ] = fresh_wire_1636[ 0 ];
	assign fresh_wire_1635[ 0 ] = fresh_wire_1594[ 0 ];
	assign fresh_wire_1637[ 0 ] = fresh_wire_1658[ 0 ];
	assign fresh_wire_1637[ 1 ] = fresh_wire_1658[ 1 ];
	assign fresh_wire_1639[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1640[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_1641[ 0 ] = fresh_wire_609[ 0 ];
	assign fresh_wire_1641[ 1 ] = fresh_wire_609[ 1 ];
	assign fresh_wire_1641[ 2 ] = fresh_wire_609[ 2 ];
	assign fresh_wire_1641[ 3 ] = fresh_wire_609[ 3 ];
	assign fresh_wire_1641[ 4 ] = fresh_wire_609[ 4 ];
	assign fresh_wire_1641[ 5 ] = fresh_wire_609[ 5 ];
	assign fresh_wire_1641[ 6 ] = fresh_wire_609[ 6 ];
	assign fresh_wire_1641[ 7 ] = fresh_wire_609[ 7 ];
	assign fresh_wire_1641[ 8 ] = fresh_wire_609[ 8 ];
	assign fresh_wire_1641[ 9 ] = fresh_wire_609[ 9 ];
	assign fresh_wire_1641[ 10 ] = fresh_wire_609[ 10 ];
	assign fresh_wire_1641[ 11 ] = fresh_wire_609[ 11 ];
	assign fresh_wire_1641[ 12 ] = fresh_wire_609[ 12 ];
	assign fresh_wire_1641[ 13 ] = fresh_wire_609[ 13 ];
	assign fresh_wire_1641[ 14 ] = fresh_wire_609[ 14 ];
	assign fresh_wire_1641[ 15 ] = fresh_wire_609[ 15 ];
	assign fresh_wire_1641[ 16 ] = fresh_wire_1642[ 0 ];
	assign fresh_wire_1641[ 17 ] = fresh_wire_1642[ 1 ];
	assign fresh_wire_1641[ 18 ] = fresh_wire_1642[ 2 ];
	assign fresh_wire_1641[ 19 ] = fresh_wire_1642[ 3 ];
	assign fresh_wire_1641[ 20 ] = fresh_wire_1642[ 4 ];
	assign fresh_wire_1641[ 21 ] = fresh_wire_1642[ 5 ];
	assign fresh_wire_1641[ 22 ] = fresh_wire_1642[ 6 ];
	assign fresh_wire_1641[ 23 ] = fresh_wire_1642[ 7 ];
	assign fresh_wire_1641[ 24 ] = fresh_wire_1642[ 8 ];
	assign fresh_wire_1641[ 25 ] = fresh_wire_1642[ 9 ];
	assign fresh_wire_1641[ 26 ] = fresh_wire_1642[ 10 ];
	assign fresh_wire_1641[ 27 ] = fresh_wire_1642[ 11 ];
	assign fresh_wire_1641[ 28 ] = fresh_wire_1642[ 12 ];
	assign fresh_wire_1641[ 29 ] = fresh_wire_1642[ 13 ];
	assign fresh_wire_1641[ 30 ] = fresh_wire_1642[ 14 ];
	assign fresh_wire_1641[ 31 ] = fresh_wire_1642[ 15 ];
	assign fresh_wire_1641[ 32 ] = fresh_wire_1642[ 16 ];
	assign fresh_wire_1641[ 33 ] = fresh_wire_1642[ 17 ];
	assign fresh_wire_1641[ 34 ] = fresh_wire_1642[ 18 ];
	assign fresh_wire_1641[ 35 ] = fresh_wire_1642[ 19 ];
	assign fresh_wire_1641[ 36 ] = fresh_wire_1642[ 20 ];
	assign fresh_wire_1641[ 37 ] = fresh_wire_1642[ 21 ];
	assign fresh_wire_1641[ 38 ] = fresh_wire_1642[ 22 ];
	assign fresh_wire_1641[ 39 ] = fresh_wire_1642[ 23 ];
	assign fresh_wire_1641[ 40 ] = fresh_wire_1642[ 24 ];
	assign fresh_wire_1641[ 41 ] = fresh_wire_1642[ 25 ];
	assign fresh_wire_1641[ 42 ] = fresh_wire_1642[ 26 ];
	assign fresh_wire_1641[ 43 ] = fresh_wire_1642[ 27 ];
	assign fresh_wire_1641[ 44 ] = fresh_wire_1642[ 28 ];
	assign fresh_wire_1641[ 45 ] = fresh_wire_1642[ 29 ];
	assign fresh_wire_1641[ 46 ] = fresh_wire_1642[ 30 ];
	assign fresh_wire_1641[ 47 ] = fresh_wire_1642[ 31 ];
	assign fresh_wire_1643[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1644[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1645[ 0 ] = fresh_wire_1597[ 0 ];
	assign fresh_wire_1647[ 0 ] = fresh_wire_1634[ 0 ];
	assign fresh_wire_1648[ 0 ] = fresh_wire_1646[ 0 ];
	assign fresh_wire_1649[ 0 ] = fresh_wire_1609[ 0 ];
	assign fresh_wire_1651[ 0 ] = fresh_wire_1629[ 0 ];
	assign fresh_wire_1652[ 0 ] = fresh_wire_1638[ 0 ];
	assign fresh_wire_1652[ 1 ] = fresh_wire_1638[ 1 ];
	assign fresh_wire_1653[ 0 ] = fresh_wire_1690[ 0 ];
	assign fresh_wire_1653[ 1 ] = fresh_wire_1690[ 1 ];
	assign fresh_wire_1655[ 0 ] = fresh_wire_1624[ 0 ];
	assign fresh_wire_1656[ 0 ] = fresh_wire_1654[ 0 ];
	assign fresh_wire_1656[ 1 ] = fresh_wire_1654[ 1 ];
	assign fresh_wire_1657[ 0 ] = fresh_wire_1585[ 0 ];
	assign fresh_wire_1657[ 1 ] = fresh_wire_1585[ 1 ];
	assign fresh_wire_1659[ 0 ] = fresh_wire_1619[ 0 ];
	assign fresh_wire_1660[ 0 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 1 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 2 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 3 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 4 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 5 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 6 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 7 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 8 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 9 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 10 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 11 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 12 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 13 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 14 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 15 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 16 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 17 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 18 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 19 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 20 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 21 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 22 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 23 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 24 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 25 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 26 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 27 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 28 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 29 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 30 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1660[ 31 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1661[ 0 ] = fresh_wire_1642[ 32 ];
	assign fresh_wire_1661[ 1 ] = fresh_wire_1642[ 33 ];
	assign fresh_wire_1661[ 2 ] = fresh_wire_1642[ 34 ];
	assign fresh_wire_1661[ 3 ] = fresh_wire_1642[ 35 ];
	assign fresh_wire_1661[ 4 ] = fresh_wire_1642[ 36 ];
	assign fresh_wire_1661[ 5 ] = fresh_wire_1642[ 37 ];
	assign fresh_wire_1661[ 6 ] = fresh_wire_1642[ 38 ];
	assign fresh_wire_1661[ 7 ] = fresh_wire_1642[ 39 ];
	assign fresh_wire_1661[ 8 ] = fresh_wire_1642[ 40 ];
	assign fresh_wire_1661[ 9 ] = fresh_wire_1642[ 41 ];
	assign fresh_wire_1661[ 10 ] = fresh_wire_1642[ 42 ];
	assign fresh_wire_1661[ 11 ] = fresh_wire_1642[ 43 ];
	assign fresh_wire_1661[ 12 ] = fresh_wire_1642[ 44 ];
	assign fresh_wire_1661[ 13 ] = fresh_wire_1642[ 45 ];
	assign fresh_wire_1661[ 14 ] = fresh_wire_1642[ 46 ];
	assign fresh_wire_1661[ 15 ] = fresh_wire_1642[ 47 ];
	assign fresh_wire_1661[ 16 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1661[ 17 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1661[ 18 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1661[ 19 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1661[ 20 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1661[ 21 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1661[ 22 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1661[ 23 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1661[ 24 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1661[ 25 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1661[ 26 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1661[ 27 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1661[ 28 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1661[ 29 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1661[ 30 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1661[ 31 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1663[ 0 ] = fresh_wire_1597[ 0 ];
	assign fresh_wire_1664[ 0 ] = fresh_wire_1662[ 0 ];
	assign fresh_wire_1664[ 1 ] = fresh_wire_1662[ 1 ];
	assign fresh_wire_1664[ 2 ] = fresh_wire_1662[ 2 ];
	assign fresh_wire_1664[ 3 ] = fresh_wire_1662[ 3 ];
	assign fresh_wire_1664[ 4 ] = fresh_wire_1662[ 4 ];
	assign fresh_wire_1664[ 5 ] = fresh_wire_1662[ 5 ];
	assign fresh_wire_1664[ 6 ] = fresh_wire_1662[ 6 ];
	assign fresh_wire_1664[ 7 ] = fresh_wire_1662[ 7 ];
	assign fresh_wire_1664[ 8 ] = fresh_wire_1662[ 8 ];
	assign fresh_wire_1664[ 9 ] = fresh_wire_1662[ 9 ];
	assign fresh_wire_1664[ 10 ] = fresh_wire_1662[ 10 ];
	assign fresh_wire_1664[ 11 ] = fresh_wire_1662[ 11 ];
	assign fresh_wire_1664[ 12 ] = fresh_wire_1662[ 12 ];
	assign fresh_wire_1664[ 13 ] = fresh_wire_1662[ 13 ];
	assign fresh_wire_1664[ 14 ] = fresh_wire_1662[ 14 ];
	assign fresh_wire_1664[ 15 ] = fresh_wire_1662[ 15 ];
	assign fresh_wire_1664[ 16 ] = fresh_wire_1662[ 16 ];
	assign fresh_wire_1664[ 17 ] = fresh_wire_1662[ 17 ];
	assign fresh_wire_1664[ 18 ] = fresh_wire_1662[ 18 ];
	assign fresh_wire_1664[ 19 ] = fresh_wire_1662[ 19 ];
	assign fresh_wire_1664[ 20 ] = fresh_wire_1662[ 20 ];
	assign fresh_wire_1664[ 21 ] = fresh_wire_1662[ 21 ];
	assign fresh_wire_1664[ 22 ] = fresh_wire_1662[ 22 ];
	assign fresh_wire_1664[ 23 ] = fresh_wire_1662[ 23 ];
	assign fresh_wire_1664[ 24 ] = fresh_wire_1662[ 24 ];
	assign fresh_wire_1664[ 25 ] = fresh_wire_1662[ 25 ];
	assign fresh_wire_1664[ 26 ] = fresh_wire_1662[ 26 ];
	assign fresh_wire_1664[ 27 ] = fresh_wire_1662[ 27 ];
	assign fresh_wire_1664[ 28 ] = fresh_wire_1662[ 28 ];
	assign fresh_wire_1664[ 29 ] = fresh_wire_1662[ 29 ];
	assign fresh_wire_1664[ 30 ] = fresh_wire_1662[ 30 ];
	assign fresh_wire_1664[ 31 ] = fresh_wire_1662[ 31 ];
	assign fresh_wire_1665[ 0 ] = fresh_wire_1642[ 16 ];
	assign fresh_wire_1665[ 1 ] = fresh_wire_1642[ 17 ];
	assign fresh_wire_1665[ 2 ] = fresh_wire_1642[ 18 ];
	assign fresh_wire_1665[ 3 ] = fresh_wire_1642[ 19 ];
	assign fresh_wire_1665[ 4 ] = fresh_wire_1642[ 20 ];
	assign fresh_wire_1665[ 5 ] = fresh_wire_1642[ 21 ];
	assign fresh_wire_1665[ 6 ] = fresh_wire_1642[ 22 ];
	assign fresh_wire_1665[ 7 ] = fresh_wire_1642[ 23 ];
	assign fresh_wire_1665[ 8 ] = fresh_wire_1642[ 24 ];
	assign fresh_wire_1665[ 9 ] = fresh_wire_1642[ 25 ];
	assign fresh_wire_1665[ 10 ] = fresh_wire_1642[ 26 ];
	assign fresh_wire_1665[ 11 ] = fresh_wire_1642[ 27 ];
	assign fresh_wire_1665[ 12 ] = fresh_wire_1642[ 28 ];
	assign fresh_wire_1665[ 13 ] = fresh_wire_1642[ 29 ];
	assign fresh_wire_1665[ 14 ] = fresh_wire_1642[ 30 ];
	assign fresh_wire_1665[ 15 ] = fresh_wire_1642[ 31 ];
	assign fresh_wire_1665[ 16 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1665[ 17 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1665[ 18 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1665[ 19 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1665[ 20 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1665[ 21 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1665[ 22 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1665[ 23 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1665[ 24 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1665[ 25 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1665[ 26 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1665[ 27 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1665[ 28 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1665[ 29 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1665[ 30 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1665[ 31 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1667[ 0 ] = fresh_wire_1600[ 0 ];
	assign fresh_wire_1668[ 0 ] = fresh_wire_1666[ 0 ];
	assign fresh_wire_1668[ 1 ] = fresh_wire_1666[ 1 ];
	assign fresh_wire_1668[ 2 ] = fresh_wire_1666[ 2 ];
	assign fresh_wire_1668[ 3 ] = fresh_wire_1666[ 3 ];
	assign fresh_wire_1668[ 4 ] = fresh_wire_1666[ 4 ];
	assign fresh_wire_1668[ 5 ] = fresh_wire_1666[ 5 ];
	assign fresh_wire_1668[ 6 ] = fresh_wire_1666[ 6 ];
	assign fresh_wire_1668[ 7 ] = fresh_wire_1666[ 7 ];
	assign fresh_wire_1668[ 8 ] = fresh_wire_1666[ 8 ];
	assign fresh_wire_1668[ 9 ] = fresh_wire_1666[ 9 ];
	assign fresh_wire_1668[ 10 ] = fresh_wire_1666[ 10 ];
	assign fresh_wire_1668[ 11 ] = fresh_wire_1666[ 11 ];
	assign fresh_wire_1668[ 12 ] = fresh_wire_1666[ 12 ];
	assign fresh_wire_1668[ 13 ] = fresh_wire_1666[ 13 ];
	assign fresh_wire_1668[ 14 ] = fresh_wire_1666[ 14 ];
	assign fresh_wire_1668[ 15 ] = fresh_wire_1666[ 15 ];
	assign fresh_wire_1668[ 16 ] = fresh_wire_1666[ 16 ];
	assign fresh_wire_1668[ 17 ] = fresh_wire_1666[ 17 ];
	assign fresh_wire_1668[ 18 ] = fresh_wire_1666[ 18 ];
	assign fresh_wire_1668[ 19 ] = fresh_wire_1666[ 19 ];
	assign fresh_wire_1668[ 20 ] = fresh_wire_1666[ 20 ];
	assign fresh_wire_1668[ 21 ] = fresh_wire_1666[ 21 ];
	assign fresh_wire_1668[ 22 ] = fresh_wire_1666[ 22 ];
	assign fresh_wire_1668[ 23 ] = fresh_wire_1666[ 23 ];
	assign fresh_wire_1668[ 24 ] = fresh_wire_1666[ 24 ];
	assign fresh_wire_1668[ 25 ] = fresh_wire_1666[ 25 ];
	assign fresh_wire_1668[ 26 ] = fresh_wire_1666[ 26 ];
	assign fresh_wire_1668[ 27 ] = fresh_wire_1666[ 27 ];
	assign fresh_wire_1668[ 28 ] = fresh_wire_1666[ 28 ];
	assign fresh_wire_1668[ 29 ] = fresh_wire_1666[ 29 ];
	assign fresh_wire_1668[ 30 ] = fresh_wire_1666[ 30 ];
	assign fresh_wire_1668[ 31 ] = fresh_wire_1666[ 31 ];
	assign fresh_wire_1669[ 0 ] = fresh_wire_1642[ 0 ];
	assign fresh_wire_1669[ 1 ] = fresh_wire_1642[ 1 ];
	assign fresh_wire_1669[ 2 ] = fresh_wire_1642[ 2 ];
	assign fresh_wire_1669[ 3 ] = fresh_wire_1642[ 3 ];
	assign fresh_wire_1669[ 4 ] = fresh_wire_1642[ 4 ];
	assign fresh_wire_1669[ 5 ] = fresh_wire_1642[ 5 ];
	assign fresh_wire_1669[ 6 ] = fresh_wire_1642[ 6 ];
	assign fresh_wire_1669[ 7 ] = fresh_wire_1642[ 7 ];
	assign fresh_wire_1669[ 8 ] = fresh_wire_1642[ 8 ];
	assign fresh_wire_1669[ 9 ] = fresh_wire_1642[ 9 ];
	assign fresh_wire_1669[ 10 ] = fresh_wire_1642[ 10 ];
	assign fresh_wire_1669[ 11 ] = fresh_wire_1642[ 11 ];
	assign fresh_wire_1669[ 12 ] = fresh_wire_1642[ 12 ];
	assign fresh_wire_1669[ 13 ] = fresh_wire_1642[ 13 ];
	assign fresh_wire_1669[ 14 ] = fresh_wire_1642[ 14 ];
	assign fresh_wire_1669[ 15 ] = fresh_wire_1642[ 15 ];
	assign fresh_wire_1669[ 16 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1669[ 17 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1669[ 18 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1669[ 19 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1669[ 20 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1669[ 21 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1669[ 22 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1669[ 23 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1669[ 24 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1669[ 25 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1669[ 26 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1669[ 27 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1669[ 28 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1669[ 29 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1669[ 30 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1669[ 31 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1671[ 0 ] = fresh_wire_1606[ 0 ];
	assign fresh_wire_1672[ 0 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 1 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 2 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 3 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 4 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 5 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 6 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 7 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 8 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 9 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 10 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 11 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 12 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 13 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 14 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 15 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 16 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 17 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 18 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 19 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 20 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 21 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 22 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 23 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 24 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 25 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 26 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 27 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 28 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 29 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 30 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1672[ 31 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1673[ 0 ] = fresh_wire_1670[ 0 ];
	assign fresh_wire_1673[ 1 ] = fresh_wire_1670[ 1 ];
	assign fresh_wire_1673[ 2 ] = fresh_wire_1670[ 2 ];
	assign fresh_wire_1673[ 3 ] = fresh_wire_1670[ 3 ];
	assign fresh_wire_1673[ 4 ] = fresh_wire_1670[ 4 ];
	assign fresh_wire_1673[ 5 ] = fresh_wire_1670[ 5 ];
	assign fresh_wire_1673[ 6 ] = fresh_wire_1670[ 6 ];
	assign fresh_wire_1673[ 7 ] = fresh_wire_1670[ 7 ];
	assign fresh_wire_1673[ 8 ] = fresh_wire_1670[ 8 ];
	assign fresh_wire_1673[ 9 ] = fresh_wire_1670[ 9 ];
	assign fresh_wire_1673[ 10 ] = fresh_wire_1670[ 10 ];
	assign fresh_wire_1673[ 11 ] = fresh_wire_1670[ 11 ];
	assign fresh_wire_1673[ 12 ] = fresh_wire_1670[ 12 ];
	assign fresh_wire_1673[ 13 ] = fresh_wire_1670[ 13 ];
	assign fresh_wire_1673[ 14 ] = fresh_wire_1670[ 14 ];
	assign fresh_wire_1673[ 15 ] = fresh_wire_1670[ 15 ];
	assign fresh_wire_1673[ 16 ] = fresh_wire_1670[ 16 ];
	assign fresh_wire_1673[ 17 ] = fresh_wire_1670[ 17 ];
	assign fresh_wire_1673[ 18 ] = fresh_wire_1670[ 18 ];
	assign fresh_wire_1673[ 19 ] = fresh_wire_1670[ 19 ];
	assign fresh_wire_1673[ 20 ] = fresh_wire_1670[ 20 ];
	assign fresh_wire_1673[ 21 ] = fresh_wire_1670[ 21 ];
	assign fresh_wire_1673[ 22 ] = fresh_wire_1670[ 22 ];
	assign fresh_wire_1673[ 23 ] = fresh_wire_1670[ 23 ];
	assign fresh_wire_1673[ 24 ] = fresh_wire_1670[ 24 ];
	assign fresh_wire_1673[ 25 ] = fresh_wire_1670[ 25 ];
	assign fresh_wire_1673[ 26 ] = fresh_wire_1670[ 26 ];
	assign fresh_wire_1673[ 27 ] = fresh_wire_1670[ 27 ];
	assign fresh_wire_1673[ 28 ] = fresh_wire_1670[ 28 ];
	assign fresh_wire_1673[ 29 ] = fresh_wire_1670[ 29 ];
	assign fresh_wire_1673[ 30 ] = fresh_wire_1670[ 30 ];
	assign fresh_wire_1673[ 31 ] = fresh_wire_1670[ 31 ];
	assign fresh_wire_1675[ 0 ] = fresh_wire_1603[ 0 ];
	assign fresh_wire_1676[ 0 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 1 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 2 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 3 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 4 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 5 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 6 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 7 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 8 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 9 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 10 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 11 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 12 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 13 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 14 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 15 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 16 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 17 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 18 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 19 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 20 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 21 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 22 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 23 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 24 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 25 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 26 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 27 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 28 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 29 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 30 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1676[ 31 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1677[ 0 ] = fresh_wire_1642[ 16 ];
	assign fresh_wire_1677[ 1 ] = fresh_wire_1642[ 17 ];
	assign fresh_wire_1677[ 2 ] = fresh_wire_1642[ 18 ];
	assign fresh_wire_1677[ 3 ] = fresh_wire_1642[ 19 ];
	assign fresh_wire_1677[ 4 ] = fresh_wire_1642[ 20 ];
	assign fresh_wire_1677[ 5 ] = fresh_wire_1642[ 21 ];
	assign fresh_wire_1677[ 6 ] = fresh_wire_1642[ 22 ];
	assign fresh_wire_1677[ 7 ] = fresh_wire_1642[ 23 ];
	assign fresh_wire_1677[ 8 ] = fresh_wire_1642[ 24 ];
	assign fresh_wire_1677[ 9 ] = fresh_wire_1642[ 25 ];
	assign fresh_wire_1677[ 10 ] = fresh_wire_1642[ 26 ];
	assign fresh_wire_1677[ 11 ] = fresh_wire_1642[ 27 ];
	assign fresh_wire_1677[ 12 ] = fresh_wire_1642[ 28 ];
	assign fresh_wire_1677[ 13 ] = fresh_wire_1642[ 29 ];
	assign fresh_wire_1677[ 14 ] = fresh_wire_1642[ 30 ];
	assign fresh_wire_1677[ 15 ] = fresh_wire_1642[ 31 ];
	assign fresh_wire_1677[ 16 ] = fresh_wire_1642[ 32 ];
	assign fresh_wire_1677[ 17 ] = fresh_wire_1642[ 33 ];
	assign fresh_wire_1677[ 18 ] = fresh_wire_1642[ 34 ];
	assign fresh_wire_1677[ 19 ] = fresh_wire_1642[ 35 ];
	assign fresh_wire_1677[ 20 ] = fresh_wire_1642[ 36 ];
	assign fresh_wire_1677[ 21 ] = fresh_wire_1642[ 37 ];
	assign fresh_wire_1677[ 22 ] = fresh_wire_1642[ 38 ];
	assign fresh_wire_1677[ 23 ] = fresh_wire_1642[ 39 ];
	assign fresh_wire_1677[ 24 ] = fresh_wire_1642[ 40 ];
	assign fresh_wire_1677[ 25 ] = fresh_wire_1642[ 41 ];
	assign fresh_wire_1677[ 26 ] = fresh_wire_1642[ 42 ];
	assign fresh_wire_1677[ 27 ] = fresh_wire_1642[ 43 ];
	assign fresh_wire_1677[ 28 ] = fresh_wire_1642[ 44 ];
	assign fresh_wire_1677[ 29 ] = fresh_wire_1642[ 45 ];
	assign fresh_wire_1677[ 30 ] = fresh_wire_1642[ 46 ];
	assign fresh_wire_1677[ 31 ] = fresh_wire_1642[ 47 ];
	assign fresh_wire_1679[ 0 ] = fresh_wire_1597[ 0 ];
	assign fresh_wire_1680[ 0 ] = fresh_wire_1678[ 0 ];
	assign fresh_wire_1680[ 1 ] = fresh_wire_1678[ 1 ];
	assign fresh_wire_1680[ 2 ] = fresh_wire_1678[ 2 ];
	assign fresh_wire_1680[ 3 ] = fresh_wire_1678[ 3 ];
	assign fresh_wire_1680[ 4 ] = fresh_wire_1678[ 4 ];
	assign fresh_wire_1680[ 5 ] = fresh_wire_1678[ 5 ];
	assign fresh_wire_1680[ 6 ] = fresh_wire_1678[ 6 ];
	assign fresh_wire_1680[ 7 ] = fresh_wire_1678[ 7 ];
	assign fresh_wire_1680[ 8 ] = fresh_wire_1678[ 8 ];
	assign fresh_wire_1680[ 9 ] = fresh_wire_1678[ 9 ];
	assign fresh_wire_1680[ 10 ] = fresh_wire_1678[ 10 ];
	assign fresh_wire_1680[ 11 ] = fresh_wire_1678[ 11 ];
	assign fresh_wire_1680[ 12 ] = fresh_wire_1678[ 12 ];
	assign fresh_wire_1680[ 13 ] = fresh_wire_1678[ 13 ];
	assign fresh_wire_1680[ 14 ] = fresh_wire_1678[ 14 ];
	assign fresh_wire_1680[ 15 ] = fresh_wire_1678[ 15 ];
	assign fresh_wire_1680[ 16 ] = fresh_wire_1678[ 16 ];
	assign fresh_wire_1680[ 17 ] = fresh_wire_1678[ 17 ];
	assign fresh_wire_1680[ 18 ] = fresh_wire_1678[ 18 ];
	assign fresh_wire_1680[ 19 ] = fresh_wire_1678[ 19 ];
	assign fresh_wire_1680[ 20 ] = fresh_wire_1678[ 20 ];
	assign fresh_wire_1680[ 21 ] = fresh_wire_1678[ 21 ];
	assign fresh_wire_1680[ 22 ] = fresh_wire_1678[ 22 ];
	assign fresh_wire_1680[ 23 ] = fresh_wire_1678[ 23 ];
	assign fresh_wire_1680[ 24 ] = fresh_wire_1678[ 24 ];
	assign fresh_wire_1680[ 25 ] = fresh_wire_1678[ 25 ];
	assign fresh_wire_1680[ 26 ] = fresh_wire_1678[ 26 ];
	assign fresh_wire_1680[ 27 ] = fresh_wire_1678[ 27 ];
	assign fresh_wire_1680[ 28 ] = fresh_wire_1678[ 28 ];
	assign fresh_wire_1680[ 29 ] = fresh_wire_1678[ 29 ];
	assign fresh_wire_1680[ 30 ] = fresh_wire_1678[ 30 ];
	assign fresh_wire_1680[ 31 ] = fresh_wire_1678[ 31 ];
	assign fresh_wire_1681[ 0 ] = fresh_wire_1642[ 0 ];
	assign fresh_wire_1681[ 1 ] = fresh_wire_1642[ 1 ];
	assign fresh_wire_1681[ 2 ] = fresh_wire_1642[ 2 ];
	assign fresh_wire_1681[ 3 ] = fresh_wire_1642[ 3 ];
	assign fresh_wire_1681[ 4 ] = fresh_wire_1642[ 4 ];
	assign fresh_wire_1681[ 5 ] = fresh_wire_1642[ 5 ];
	assign fresh_wire_1681[ 6 ] = fresh_wire_1642[ 6 ];
	assign fresh_wire_1681[ 7 ] = fresh_wire_1642[ 7 ];
	assign fresh_wire_1681[ 8 ] = fresh_wire_1642[ 8 ];
	assign fresh_wire_1681[ 9 ] = fresh_wire_1642[ 9 ];
	assign fresh_wire_1681[ 10 ] = fresh_wire_1642[ 10 ];
	assign fresh_wire_1681[ 11 ] = fresh_wire_1642[ 11 ];
	assign fresh_wire_1681[ 12 ] = fresh_wire_1642[ 12 ];
	assign fresh_wire_1681[ 13 ] = fresh_wire_1642[ 13 ];
	assign fresh_wire_1681[ 14 ] = fresh_wire_1642[ 14 ];
	assign fresh_wire_1681[ 15 ] = fresh_wire_1642[ 15 ];
	assign fresh_wire_1681[ 16 ] = fresh_wire_1642[ 16 ];
	assign fresh_wire_1681[ 17 ] = fresh_wire_1642[ 17 ];
	assign fresh_wire_1681[ 18 ] = fresh_wire_1642[ 18 ];
	assign fresh_wire_1681[ 19 ] = fresh_wire_1642[ 19 ];
	assign fresh_wire_1681[ 20 ] = fresh_wire_1642[ 20 ];
	assign fresh_wire_1681[ 21 ] = fresh_wire_1642[ 21 ];
	assign fresh_wire_1681[ 22 ] = fresh_wire_1642[ 22 ];
	assign fresh_wire_1681[ 23 ] = fresh_wire_1642[ 23 ];
	assign fresh_wire_1681[ 24 ] = fresh_wire_1642[ 24 ];
	assign fresh_wire_1681[ 25 ] = fresh_wire_1642[ 25 ];
	assign fresh_wire_1681[ 26 ] = fresh_wire_1642[ 26 ];
	assign fresh_wire_1681[ 27 ] = fresh_wire_1642[ 27 ];
	assign fresh_wire_1681[ 28 ] = fresh_wire_1642[ 28 ];
	assign fresh_wire_1681[ 29 ] = fresh_wire_1642[ 29 ];
	assign fresh_wire_1681[ 30 ] = fresh_wire_1642[ 30 ];
	assign fresh_wire_1681[ 31 ] = fresh_wire_1642[ 31 ];
	assign fresh_wire_1683[ 0 ] = fresh_wire_1600[ 0 ];
	assign fresh_wire_1684[ 0 ] = fresh_wire_1674[ 0 ];
	assign fresh_wire_1684[ 1 ] = fresh_wire_1674[ 1 ];
	assign fresh_wire_1684[ 2 ] = fresh_wire_1674[ 2 ];
	assign fresh_wire_1684[ 3 ] = fresh_wire_1674[ 3 ];
	assign fresh_wire_1684[ 4 ] = fresh_wire_1674[ 4 ];
	assign fresh_wire_1684[ 5 ] = fresh_wire_1674[ 5 ];
	assign fresh_wire_1684[ 6 ] = fresh_wire_1674[ 6 ];
	assign fresh_wire_1684[ 7 ] = fresh_wire_1674[ 7 ];
	assign fresh_wire_1684[ 8 ] = fresh_wire_1674[ 8 ];
	assign fresh_wire_1684[ 9 ] = fresh_wire_1674[ 9 ];
	assign fresh_wire_1684[ 10 ] = fresh_wire_1674[ 10 ];
	assign fresh_wire_1684[ 11 ] = fresh_wire_1674[ 11 ];
	assign fresh_wire_1684[ 12 ] = fresh_wire_1674[ 12 ];
	assign fresh_wire_1684[ 13 ] = fresh_wire_1674[ 13 ];
	assign fresh_wire_1684[ 14 ] = fresh_wire_1674[ 14 ];
	assign fresh_wire_1684[ 15 ] = fresh_wire_1674[ 15 ];
	assign fresh_wire_1684[ 16 ] = fresh_wire_1674[ 16 ];
	assign fresh_wire_1684[ 17 ] = fresh_wire_1674[ 17 ];
	assign fresh_wire_1684[ 18 ] = fresh_wire_1674[ 18 ];
	assign fresh_wire_1684[ 19 ] = fresh_wire_1674[ 19 ];
	assign fresh_wire_1684[ 20 ] = fresh_wire_1674[ 20 ];
	assign fresh_wire_1684[ 21 ] = fresh_wire_1674[ 21 ];
	assign fresh_wire_1684[ 22 ] = fresh_wire_1674[ 22 ];
	assign fresh_wire_1684[ 23 ] = fresh_wire_1674[ 23 ];
	assign fresh_wire_1684[ 24 ] = fresh_wire_1674[ 24 ];
	assign fresh_wire_1684[ 25 ] = fresh_wire_1674[ 25 ];
	assign fresh_wire_1684[ 26 ] = fresh_wire_1674[ 26 ];
	assign fresh_wire_1684[ 27 ] = fresh_wire_1674[ 27 ];
	assign fresh_wire_1684[ 28 ] = fresh_wire_1674[ 28 ];
	assign fresh_wire_1684[ 29 ] = fresh_wire_1674[ 29 ];
	assign fresh_wire_1684[ 30 ] = fresh_wire_1674[ 30 ];
	assign fresh_wire_1684[ 31 ] = fresh_wire_1674[ 31 ];
	assign fresh_wire_1685[ 0 ] = fresh_wire_1682[ 0 ];
	assign fresh_wire_1685[ 1 ] = fresh_wire_1682[ 1 ];
	assign fresh_wire_1685[ 2 ] = fresh_wire_1682[ 2 ];
	assign fresh_wire_1685[ 3 ] = fresh_wire_1682[ 3 ];
	assign fresh_wire_1685[ 4 ] = fresh_wire_1682[ 4 ];
	assign fresh_wire_1685[ 5 ] = fresh_wire_1682[ 5 ];
	assign fresh_wire_1685[ 6 ] = fresh_wire_1682[ 6 ];
	assign fresh_wire_1685[ 7 ] = fresh_wire_1682[ 7 ];
	assign fresh_wire_1685[ 8 ] = fresh_wire_1682[ 8 ];
	assign fresh_wire_1685[ 9 ] = fresh_wire_1682[ 9 ];
	assign fresh_wire_1685[ 10 ] = fresh_wire_1682[ 10 ];
	assign fresh_wire_1685[ 11 ] = fresh_wire_1682[ 11 ];
	assign fresh_wire_1685[ 12 ] = fresh_wire_1682[ 12 ];
	assign fresh_wire_1685[ 13 ] = fresh_wire_1682[ 13 ];
	assign fresh_wire_1685[ 14 ] = fresh_wire_1682[ 14 ];
	assign fresh_wire_1685[ 15 ] = fresh_wire_1682[ 15 ];
	assign fresh_wire_1685[ 16 ] = fresh_wire_1682[ 16 ];
	assign fresh_wire_1685[ 17 ] = fresh_wire_1682[ 17 ];
	assign fresh_wire_1685[ 18 ] = fresh_wire_1682[ 18 ];
	assign fresh_wire_1685[ 19 ] = fresh_wire_1682[ 19 ];
	assign fresh_wire_1685[ 20 ] = fresh_wire_1682[ 20 ];
	assign fresh_wire_1685[ 21 ] = fresh_wire_1682[ 21 ];
	assign fresh_wire_1685[ 22 ] = fresh_wire_1682[ 22 ];
	assign fresh_wire_1685[ 23 ] = fresh_wire_1682[ 23 ];
	assign fresh_wire_1685[ 24 ] = fresh_wire_1682[ 24 ];
	assign fresh_wire_1685[ 25 ] = fresh_wire_1682[ 25 ];
	assign fresh_wire_1685[ 26 ] = fresh_wire_1682[ 26 ];
	assign fresh_wire_1685[ 27 ] = fresh_wire_1682[ 27 ];
	assign fresh_wire_1685[ 28 ] = fresh_wire_1682[ 28 ];
	assign fresh_wire_1685[ 29 ] = fresh_wire_1682[ 29 ];
	assign fresh_wire_1685[ 30 ] = fresh_wire_1682[ 30 ];
	assign fresh_wire_1685[ 31 ] = fresh_wire_1682[ 31 ];
	assign fresh_wire_1687[ 0 ] = fresh_wire_1594[ 0 ];
	assign fresh_wire_1688[ 0 ] = fresh_wire_1638[ 0 ];
	assign fresh_wire_1688[ 1 ] = fresh_wire_1638[ 1 ];
	assign fresh_wire_1689[ 0 ] = fresh_wire_1691[ 0 ];
	assign fresh_wire_1689[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1692[ 0 ] = fresh_wire_1830[ 0 ];
	assign fresh_wire_1692[ 1 ] = fresh_wire_1830[ 1 ];
	assign fresh_wire_1693[ 0 ] = fresh_wire_1899[ 0 ];
	assign fresh_wire_1693[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1695[ 0 ] = fresh_wire_1830[ 0 ];
	assign fresh_wire_1695[ 1 ] = fresh_wire_1830[ 1 ];
	assign fresh_wire_1696[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1696[ 1 ] = fresh_wire_1899[ 0 ];
	assign fresh_wire_1698[ 0 ] = fresh_wire_1358[ 0 ];
	assign fresh_wire_1699[ 0 ] = fresh_wire_1899[ 0 ];
	assign fresh_wire_1701[ 0 ] = fresh_wire_1354[ 0 ];
	assign fresh_wire_1702[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1704[ 0 ] = fresh_wire_1362[ 0 ];
	assign fresh_wire_1705[ 0 ] = fresh_wire_1899[ 0 ];
	assign fresh_wire_1707[ 0 ] = fresh_wire_1354[ 0 ];
	assign fresh_wire_1708[ 0 ] = fresh_wire_1899[ 0 ];
	assign fresh_wire_1710[ 0 ] = fresh_wire_1358[ 0 ];
	assign fresh_wire_1711[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1713[ 0 ] = fresh_wire_1362[ 0 ];
	assign fresh_wire_1714[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1716[ 0 ] = fresh_wire_1830[ 0 ];
	assign fresh_wire_1716[ 1 ] = fresh_wire_1830[ 1 ];
	assign fresh_wire_1717[ 0 ] = fresh_wire_1899[ 0 ];
	assign fresh_wire_1717[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1719[ 0 ] = fresh_wire_1830[ 0 ];
	assign fresh_wire_1719[ 1 ] = fresh_wire_1830[ 1 ];
	assign fresh_wire_1720[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1720[ 1 ] = fresh_wire_1899[ 0 ];
	assign fresh_wire_1722[ 0 ] = fresh_wire_1830[ 0 ];
	assign fresh_wire_1722[ 1 ] = fresh_wire_1830[ 1 ];
	assign fresh_wire_1723[ 0 ] = fresh_wire_1899[ 0 ];
	assign fresh_wire_1723[ 1 ] = fresh_wire_1899[ 0 ];
	assign fresh_wire_1725[ 0 ] = fresh_wire_1830[ 0 ];
	assign fresh_wire_1725[ 1 ] = fresh_wire_1830[ 1 ];
	assign fresh_wire_1726[ 0 ] = fresh_wire_1899[ 0 ];
	assign fresh_wire_1726[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1728[ 0 ] = fresh_wire_1830[ 0 ];
	assign fresh_wire_1728[ 1 ] = fresh_wire_1830[ 1 ];
	assign fresh_wire_1729[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1729[ 1 ] = fresh_wire_1899[ 0 ];
	assign fresh_wire_1731[ 0 ] = fresh_wire_1700[ 0 ];
	assign fresh_wire_1733[ 0 ] = fresh_wire_1732[ 0 ];
	assign fresh_wire_1734[ 0 ] = fresh_wire_1737[ 0 ];
	assign fresh_wire_1736[ 0 ] = fresh_wire_1703[ 0 ];
	assign fresh_wire_1738[ 0 ] = fresh_wire_1706[ 0 ];
	assign fresh_wire_1740[ 0 ] = fresh_wire_1739[ 0 ];
	assign fresh_wire_1741[ 0 ] = fresh_wire_1744[ 0 ];
	assign fresh_wire_1743[ 0 ] = fresh_wire_1703[ 0 ];
	assign fresh_wire_1745[ 0 ] = fresh_wire_1700[ 0 ];
	assign fresh_wire_1747[ 0 ] = fresh_wire_1746[ 0 ];
	assign fresh_wire_1748[ 0 ] = fresh_wire_1751[ 0 ];
	assign fresh_wire_1750[ 0 ] = fresh_wire_1709[ 0 ];
	assign fresh_wire_1752[ 0 ] = fresh_wire_1706[ 0 ];
	assign fresh_wire_1754[ 0 ] = fresh_wire_1753[ 0 ];
	assign fresh_wire_1755[ 0 ] = fresh_wire_1758[ 0 ];
	assign fresh_wire_1757[ 0 ] = fresh_wire_1709[ 0 ];
	assign fresh_wire_1759[ 0 ] = fresh_wire_1712[ 0 ];
	assign fresh_wire_1761[ 0 ] = fresh_wire_1760[ 0 ];
	assign fresh_wire_1762[ 0 ] = fresh_wire_1765[ 0 ];
	assign fresh_wire_1764[ 0 ] = fresh_wire_1715[ 0 ];
	assign fresh_wire_1766[ 0 ] = fresh_wire_1763[ 0 ];
	assign fresh_wire_1768[ 0 ] = fresh_wire_1767[ 0 ];
	assign fresh_wire_1769[ 0 ] = fresh_wire_1772[ 0 ];
	assign fresh_wire_1771[ 0 ] = fresh_wire_1703[ 0 ];
	assign fresh_wire_1773[ 0 ] = fresh_wire_1712[ 0 ];
	assign fresh_wire_1775[ 0 ] = fresh_wire_1774[ 0 ];
	assign fresh_wire_1776[ 0 ] = fresh_wire_1779[ 0 ];
	assign fresh_wire_1778[ 0 ] = fresh_wire_1715[ 0 ];
	assign fresh_wire_1780[ 0 ] = fresh_wire_1777[ 0 ];
	assign fresh_wire_1782[ 0 ] = fresh_wire_1781[ 0 ];
	assign fresh_wire_1783[ 0 ] = fresh_wire_1786[ 0 ];
	assign fresh_wire_1785[ 0 ] = fresh_wire_1709[ 0 ];
	assign fresh_wire_1787[ 0 ] = fresh_wire_1821[ 0 ];
	assign fresh_wire_1789[ 0 ] = fresh_wire_1788[ 0 ];
	assign fresh_wire_1790[ 0 ] = fresh_wire_1793[ 0 ];
	assign fresh_wire_1792[ 0 ] = fresh_wire_1703[ 0 ];
	assign fresh_wire_1794[ 0 ] = fresh_wire_1828[ 0 ];
	assign fresh_wire_1796[ 0 ] = fresh_wire_1795[ 0 ];
	assign fresh_wire_1797[ 0 ] = fresh_wire_1800[ 0 ];
	assign fresh_wire_1799[ 0 ] = fresh_wire_1709[ 0 ];
	assign fresh_wire_1801[ 0 ] = fresh_wire_1712[ 0 ];
	assign fresh_wire_1803[ 0 ] = fresh_wire_1802[ 0 ];
	assign fresh_wire_1804[ 0 ] = fresh_wire_1807[ 0 ];
	assign fresh_wire_1806[ 0 ] = fresh_wire_1715[ 0 ];
	assign fresh_wire_1808[ 0 ] = fresh_wire_1805[ 0 ];
	assign fresh_wire_1810[ 0 ] = fresh_wire_1809[ 0 ];
	assign fresh_wire_1811[ 0 ] = fresh_wire_1814[ 0 ];
	assign fresh_wire_1813[ 0 ] = fresh_wire_1709[ 0 ];
	assign fresh_wire_1815[ 0 ] = fresh_wire_1700[ 0 ];
	assign fresh_wire_1817[ 0 ] = fresh_wire_1706[ 0 ];
	assign fresh_wire_1819[ 0 ] = fresh_wire_1816[ 0 ];
	assign fresh_wire_1820[ 0 ] = fresh_wire_1818[ 0 ];
	assign fresh_wire_1822[ 0 ] = fresh_wire_1700[ 0 ];
	assign fresh_wire_1824[ 0 ] = fresh_wire_1706[ 0 ];
	assign fresh_wire_1826[ 0 ] = fresh_wire_1823[ 0 ];
	assign fresh_wire_1827[ 0 ] = fresh_wire_1825[ 0 ];
	assign fresh_wire_1829[ 0 ] = fresh_wire_1886[ 0 ];
	assign fresh_wire_1829[ 1 ] = fresh_wire_1886[ 1 ];
	assign fresh_wire_1831[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1832[ 0 ] = fresh_wire_2250[ 0 ];
	assign fresh_wire_1833[ 0 ] = fresh_wire_1894[ 0 ];
	assign fresh_wire_1833[ 1 ] = fresh_wire_1894[ 1 ];
	assign fresh_wire_1833[ 2 ] = fresh_wire_1894[ 2 ];
	assign fresh_wire_1833[ 3 ] = fresh_wire_1894[ 3 ];
	assign fresh_wire_1833[ 4 ] = fresh_wire_1894[ 4 ];
	assign fresh_wire_1833[ 5 ] = fresh_wire_1894[ 5 ];
	assign fresh_wire_1833[ 6 ] = fresh_wire_1894[ 6 ];
	assign fresh_wire_1833[ 7 ] = fresh_wire_1894[ 7 ];
	assign fresh_wire_1833[ 8 ] = fresh_wire_1894[ 8 ];
	assign fresh_wire_1833[ 9 ] = fresh_wire_1894[ 9 ];
	assign fresh_wire_1833[ 10 ] = fresh_wire_1894[ 10 ];
	assign fresh_wire_1833[ 11 ] = fresh_wire_1894[ 11 ];
	assign fresh_wire_1833[ 12 ] = fresh_wire_1894[ 12 ];
	assign fresh_wire_1833[ 13 ] = fresh_wire_1894[ 13 ];
	assign fresh_wire_1833[ 14 ] = fresh_wire_1894[ 14 ];
	assign fresh_wire_1833[ 15 ] = fresh_wire_1894[ 15 ];
	assign fresh_wire_1833[ 16 ] = fresh_wire_1894[ 16 ];
	assign fresh_wire_1833[ 17 ] = fresh_wire_1894[ 17 ];
	assign fresh_wire_1833[ 18 ] = fresh_wire_1894[ 18 ];
	assign fresh_wire_1833[ 19 ] = fresh_wire_1894[ 19 ];
	assign fresh_wire_1833[ 20 ] = fresh_wire_1894[ 20 ];
	assign fresh_wire_1833[ 21 ] = fresh_wire_1894[ 21 ];
	assign fresh_wire_1833[ 22 ] = fresh_wire_1894[ 22 ];
	assign fresh_wire_1833[ 23 ] = fresh_wire_1894[ 23 ];
	assign fresh_wire_1833[ 24 ] = fresh_wire_1894[ 24 ];
	assign fresh_wire_1833[ 25 ] = fresh_wire_1894[ 25 ];
	assign fresh_wire_1833[ 26 ] = fresh_wire_1894[ 26 ];
	assign fresh_wire_1833[ 27 ] = fresh_wire_1894[ 27 ];
	assign fresh_wire_1833[ 28 ] = fresh_wire_1894[ 28 ];
	assign fresh_wire_1833[ 29 ] = fresh_wire_1894[ 29 ];
	assign fresh_wire_1833[ 30 ] = fresh_wire_1894[ 30 ];
	assign fresh_wire_1833[ 31 ] = fresh_wire_1894[ 31 ];
	assign fresh_wire_1833[ 32 ] = fresh_wire_1894[ 32 ];
	assign fresh_wire_1833[ 33 ] = fresh_wire_1894[ 33 ];
	assign fresh_wire_1833[ 34 ] = fresh_wire_1894[ 34 ];
	assign fresh_wire_1833[ 35 ] = fresh_wire_1894[ 35 ];
	assign fresh_wire_1833[ 36 ] = fresh_wire_1894[ 36 ];
	assign fresh_wire_1833[ 37 ] = fresh_wire_1894[ 37 ];
	assign fresh_wire_1833[ 38 ] = fresh_wire_1894[ 38 ];
	assign fresh_wire_1833[ 39 ] = fresh_wire_1894[ 39 ];
	assign fresh_wire_1833[ 40 ] = fresh_wire_1894[ 40 ];
	assign fresh_wire_1833[ 41 ] = fresh_wire_1894[ 41 ];
	assign fresh_wire_1833[ 42 ] = fresh_wire_1894[ 42 ];
	assign fresh_wire_1833[ 43 ] = fresh_wire_1894[ 43 ];
	assign fresh_wire_1833[ 44 ] = fresh_wire_1894[ 44 ];
	assign fresh_wire_1833[ 45 ] = fresh_wire_1894[ 45 ];
	assign fresh_wire_1833[ 46 ] = fresh_wire_1894[ 46 ];
	assign fresh_wire_1833[ 47 ] = fresh_wire_1894[ 47 ];
	assign fresh_wire_1835[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1836[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1836[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1836[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1836[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1836[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1836[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1836[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1836[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1836[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1836[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1836[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1836[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1836[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1836[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1836[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1836[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1837[ 0 ] = fresh_wire_1834[ 32 ];
	assign fresh_wire_1837[ 1 ] = fresh_wire_1834[ 33 ];
	assign fresh_wire_1837[ 2 ] = fresh_wire_1834[ 34 ];
	assign fresh_wire_1837[ 3 ] = fresh_wire_1834[ 35 ];
	assign fresh_wire_1837[ 4 ] = fresh_wire_1834[ 36 ];
	assign fresh_wire_1837[ 5 ] = fresh_wire_1834[ 37 ];
	assign fresh_wire_1837[ 6 ] = fresh_wire_1834[ 38 ];
	assign fresh_wire_1837[ 7 ] = fresh_wire_1834[ 39 ];
	assign fresh_wire_1837[ 8 ] = fresh_wire_1834[ 40 ];
	assign fresh_wire_1837[ 9 ] = fresh_wire_1834[ 41 ];
	assign fresh_wire_1837[ 10 ] = fresh_wire_1834[ 42 ];
	assign fresh_wire_1837[ 11 ] = fresh_wire_1834[ 43 ];
	assign fresh_wire_1837[ 12 ] = fresh_wire_1834[ 44 ];
	assign fresh_wire_1837[ 13 ] = fresh_wire_1834[ 45 ];
	assign fresh_wire_1837[ 14 ] = fresh_wire_1834[ 46 ];
	assign fresh_wire_1837[ 15 ] = fresh_wire_1834[ 47 ];
	assign fresh_wire_1839[ 0 ] = fresh_wire_1724[ 0 ];
	assign fresh_wire_1840[ 0 ] = fresh_wire_1838[ 0 ];
	assign fresh_wire_1840[ 1 ] = fresh_wire_1838[ 1 ];
	assign fresh_wire_1840[ 2 ] = fresh_wire_1838[ 2 ];
	assign fresh_wire_1840[ 3 ] = fresh_wire_1838[ 3 ];
	assign fresh_wire_1840[ 4 ] = fresh_wire_1838[ 4 ];
	assign fresh_wire_1840[ 5 ] = fresh_wire_1838[ 5 ];
	assign fresh_wire_1840[ 6 ] = fresh_wire_1838[ 6 ];
	assign fresh_wire_1840[ 7 ] = fresh_wire_1838[ 7 ];
	assign fresh_wire_1840[ 8 ] = fresh_wire_1838[ 8 ];
	assign fresh_wire_1840[ 9 ] = fresh_wire_1838[ 9 ];
	assign fresh_wire_1840[ 10 ] = fresh_wire_1838[ 10 ];
	assign fresh_wire_1840[ 11 ] = fresh_wire_1838[ 11 ];
	assign fresh_wire_1840[ 12 ] = fresh_wire_1838[ 12 ];
	assign fresh_wire_1840[ 13 ] = fresh_wire_1838[ 13 ];
	assign fresh_wire_1840[ 14 ] = fresh_wire_1838[ 14 ];
	assign fresh_wire_1840[ 15 ] = fresh_wire_1838[ 15 ];
	assign fresh_wire_1841[ 0 ] = fresh_wire_1834[ 16 ];
	assign fresh_wire_1841[ 1 ] = fresh_wire_1834[ 17 ];
	assign fresh_wire_1841[ 2 ] = fresh_wire_1834[ 18 ];
	assign fresh_wire_1841[ 3 ] = fresh_wire_1834[ 19 ];
	assign fresh_wire_1841[ 4 ] = fresh_wire_1834[ 20 ];
	assign fresh_wire_1841[ 5 ] = fresh_wire_1834[ 21 ];
	assign fresh_wire_1841[ 6 ] = fresh_wire_1834[ 22 ];
	assign fresh_wire_1841[ 7 ] = fresh_wire_1834[ 23 ];
	assign fresh_wire_1841[ 8 ] = fresh_wire_1834[ 24 ];
	assign fresh_wire_1841[ 9 ] = fresh_wire_1834[ 25 ];
	assign fresh_wire_1841[ 10 ] = fresh_wire_1834[ 26 ];
	assign fresh_wire_1841[ 11 ] = fresh_wire_1834[ 27 ];
	assign fresh_wire_1841[ 12 ] = fresh_wire_1834[ 28 ];
	assign fresh_wire_1841[ 13 ] = fresh_wire_1834[ 29 ];
	assign fresh_wire_1841[ 14 ] = fresh_wire_1834[ 30 ];
	assign fresh_wire_1841[ 15 ] = fresh_wire_1834[ 31 ];
	assign fresh_wire_1843[ 0 ] = fresh_wire_1721[ 0 ];
	assign fresh_wire_1844[ 0 ] = fresh_wire_1842[ 0 ];
	assign fresh_wire_1844[ 1 ] = fresh_wire_1842[ 1 ];
	assign fresh_wire_1844[ 2 ] = fresh_wire_1842[ 2 ];
	assign fresh_wire_1844[ 3 ] = fresh_wire_1842[ 3 ];
	assign fresh_wire_1844[ 4 ] = fresh_wire_1842[ 4 ];
	assign fresh_wire_1844[ 5 ] = fresh_wire_1842[ 5 ];
	assign fresh_wire_1844[ 6 ] = fresh_wire_1842[ 6 ];
	assign fresh_wire_1844[ 7 ] = fresh_wire_1842[ 7 ];
	assign fresh_wire_1844[ 8 ] = fresh_wire_1842[ 8 ];
	assign fresh_wire_1844[ 9 ] = fresh_wire_1842[ 9 ];
	assign fresh_wire_1844[ 10 ] = fresh_wire_1842[ 10 ];
	assign fresh_wire_1844[ 11 ] = fresh_wire_1842[ 11 ];
	assign fresh_wire_1844[ 12 ] = fresh_wire_1842[ 12 ];
	assign fresh_wire_1844[ 13 ] = fresh_wire_1842[ 13 ];
	assign fresh_wire_1844[ 14 ] = fresh_wire_1842[ 14 ];
	assign fresh_wire_1844[ 15 ] = fresh_wire_1842[ 15 ];
	assign fresh_wire_1845[ 0 ] = fresh_wire_1834[ 0 ];
	assign fresh_wire_1845[ 1 ] = fresh_wire_1834[ 1 ];
	assign fresh_wire_1845[ 2 ] = fresh_wire_1834[ 2 ];
	assign fresh_wire_1845[ 3 ] = fresh_wire_1834[ 3 ];
	assign fresh_wire_1845[ 4 ] = fresh_wire_1834[ 4 ];
	assign fresh_wire_1845[ 5 ] = fresh_wire_1834[ 5 ];
	assign fresh_wire_1845[ 6 ] = fresh_wire_1834[ 6 ];
	assign fresh_wire_1845[ 7 ] = fresh_wire_1834[ 7 ];
	assign fresh_wire_1845[ 8 ] = fresh_wire_1834[ 8 ];
	assign fresh_wire_1845[ 9 ] = fresh_wire_1834[ 9 ];
	assign fresh_wire_1845[ 10 ] = fresh_wire_1834[ 10 ];
	assign fresh_wire_1845[ 11 ] = fresh_wire_1834[ 11 ];
	assign fresh_wire_1845[ 12 ] = fresh_wire_1834[ 12 ];
	assign fresh_wire_1845[ 13 ] = fresh_wire_1834[ 13 ];
	assign fresh_wire_1845[ 14 ] = fresh_wire_1834[ 14 ];
	assign fresh_wire_1845[ 15 ] = fresh_wire_1834[ 15 ];
	assign fresh_wire_1847[ 0 ] = fresh_wire_1718[ 0 ];
	assign fresh_wire_1848[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1848[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1848[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1848[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1848[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1848[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1848[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1848[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1848[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1848[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1848[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1848[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1848[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1848[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1848[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1848[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1849[ 0 ] = fresh_wire_1846[ 0 ];
	assign fresh_wire_1849[ 1 ] = fresh_wire_1846[ 1 ];
	assign fresh_wire_1849[ 2 ] = fresh_wire_1846[ 2 ];
	assign fresh_wire_1849[ 3 ] = fresh_wire_1846[ 3 ];
	assign fresh_wire_1849[ 4 ] = fresh_wire_1846[ 4 ];
	assign fresh_wire_1849[ 5 ] = fresh_wire_1846[ 5 ];
	assign fresh_wire_1849[ 6 ] = fresh_wire_1846[ 6 ];
	assign fresh_wire_1849[ 7 ] = fresh_wire_1846[ 7 ];
	assign fresh_wire_1849[ 8 ] = fresh_wire_1846[ 8 ];
	assign fresh_wire_1849[ 9 ] = fresh_wire_1846[ 9 ];
	assign fresh_wire_1849[ 10 ] = fresh_wire_1846[ 10 ];
	assign fresh_wire_1849[ 11 ] = fresh_wire_1846[ 11 ];
	assign fresh_wire_1849[ 12 ] = fresh_wire_1846[ 12 ];
	assign fresh_wire_1849[ 13 ] = fresh_wire_1846[ 13 ];
	assign fresh_wire_1849[ 14 ] = fresh_wire_1846[ 14 ];
	assign fresh_wire_1849[ 15 ] = fresh_wire_1846[ 15 ];
	assign fresh_wire_1851[ 0 ] = fresh_wire_1709[ 0 ];
	assign fresh_wire_1852[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1853[ 0 ] = fresh_wire_1899[ 0 ];
	assign fresh_wire_1855[ 0 ] = fresh_wire_1798[ 0 ];
	assign fresh_wire_1856[ 0 ] = fresh_wire_1854[ 0 ];
	assign fresh_wire_1857[ 0 ] = fresh_wire_1899[ 0 ];
	assign fresh_wire_1859[ 0 ] = fresh_wire_1791[ 0 ];
	assign fresh_wire_1860[ 0 ] = fresh_wire_1858[ 0 ];
	assign fresh_wire_1861[ 0 ] = fresh_wire_1730[ 0 ];
	assign fresh_wire_1863[ 0 ] = fresh_wire_1784[ 0 ];
	assign fresh_wire_1864[ 0 ] = fresh_wire_1862[ 0 ];
	assign fresh_wire_1865[ 0 ] = fresh_wire_1727[ 0 ];
	assign fresh_wire_1867[ 0 ] = fresh_wire_1770[ 0 ];
	assign fresh_wire_1868[ 0 ] = fresh_wire_1830[ 0 ];
	assign fresh_wire_1868[ 1 ] = fresh_wire_1830[ 1 ];
	assign fresh_wire_1869[ 0 ] = fresh_wire_1694[ 0 ];
	assign fresh_wire_1869[ 1 ] = fresh_wire_1694[ 1 ];
	assign fresh_wire_1871[ 0 ] = fresh_wire_1756[ 0 ];
	assign fresh_wire_1872[ 0 ] = fresh_wire_1870[ 0 ];
	assign fresh_wire_1872[ 1 ] = fresh_wire_1870[ 1 ];
	assign fresh_wire_1873[ 0 ] = fresh_wire_1830[ 0 ];
	assign fresh_wire_1873[ 1 ] = fresh_wire_1830[ 1 ];
	assign fresh_wire_1875[ 0 ] = fresh_wire_1749[ 0 ];
	assign fresh_wire_1876[ 0 ] = fresh_wire_1874[ 0 ];
	assign fresh_wire_1876[ 1 ] = fresh_wire_1874[ 1 ];
	assign fresh_wire_1877[ 0 ] = fresh_wire_1697[ 0 ];
	assign fresh_wire_1877[ 1 ] = fresh_wire_1697[ 1 ];
	assign fresh_wire_1879[ 0 ] = fresh_wire_1742[ 0 ];
	assign fresh_wire_1880[ 0 ] = fresh_wire_1878[ 0 ];
	assign fresh_wire_1880[ 1 ] = fresh_wire_1878[ 1 ];
	assign fresh_wire_1881[ 0 ] = fresh_wire_1694[ 0 ];
	assign fresh_wire_1881[ 1 ] = fresh_wire_1694[ 1 ];
	assign fresh_wire_1883[ 0 ] = fresh_wire_1735[ 0 ];
	assign fresh_wire_1884[ 0 ] = fresh_wire_1882[ 0 ];
	assign fresh_wire_1884[ 1 ] = fresh_wire_1882[ 1 ];
	assign fresh_wire_1885[ 0 ] = fresh_wire_1898[ 0 ];
	assign fresh_wire_1885[ 1 ] = fresh_wire_1898[ 1 ];
	assign fresh_wire_1887[ 0 ] = fresh_wire_1812[ 0 ];
	assign fresh_wire_1888[ 0 ] = fresh_wire_1834[ 0 ];
	assign fresh_wire_1888[ 1 ] = fresh_wire_1834[ 1 ];
	assign fresh_wire_1888[ 2 ] = fresh_wire_1834[ 2 ];
	assign fresh_wire_1888[ 3 ] = fresh_wire_1834[ 3 ];
	assign fresh_wire_1888[ 4 ] = fresh_wire_1834[ 4 ];
	assign fresh_wire_1888[ 5 ] = fresh_wire_1834[ 5 ];
	assign fresh_wire_1888[ 6 ] = fresh_wire_1834[ 6 ];
	assign fresh_wire_1888[ 7 ] = fresh_wire_1834[ 7 ];
	assign fresh_wire_1888[ 8 ] = fresh_wire_1834[ 8 ];
	assign fresh_wire_1888[ 9 ] = fresh_wire_1834[ 9 ];
	assign fresh_wire_1888[ 10 ] = fresh_wire_1834[ 10 ];
	assign fresh_wire_1888[ 11 ] = fresh_wire_1834[ 11 ];
	assign fresh_wire_1888[ 12 ] = fresh_wire_1834[ 12 ];
	assign fresh_wire_1888[ 13 ] = fresh_wire_1834[ 13 ];
	assign fresh_wire_1888[ 14 ] = fresh_wire_1834[ 14 ];
	assign fresh_wire_1888[ 15 ] = fresh_wire_1834[ 15 ];
	assign fresh_wire_1888[ 16 ] = fresh_wire_1834[ 16 ];
	assign fresh_wire_1888[ 17 ] = fresh_wire_1834[ 17 ];
	assign fresh_wire_1888[ 18 ] = fresh_wire_1834[ 18 ];
	assign fresh_wire_1888[ 19 ] = fresh_wire_1834[ 19 ];
	assign fresh_wire_1888[ 20 ] = fresh_wire_1834[ 20 ];
	assign fresh_wire_1888[ 21 ] = fresh_wire_1834[ 21 ];
	assign fresh_wire_1888[ 22 ] = fresh_wire_1834[ 22 ];
	assign fresh_wire_1888[ 23 ] = fresh_wire_1834[ 23 ];
	assign fresh_wire_1888[ 24 ] = fresh_wire_1834[ 24 ];
	assign fresh_wire_1888[ 25 ] = fresh_wire_1834[ 25 ];
	assign fresh_wire_1888[ 26 ] = fresh_wire_1834[ 26 ];
	assign fresh_wire_1888[ 27 ] = fresh_wire_1834[ 27 ];
	assign fresh_wire_1888[ 28 ] = fresh_wire_1834[ 28 ];
	assign fresh_wire_1888[ 29 ] = fresh_wire_1834[ 29 ];
	assign fresh_wire_1888[ 30 ] = fresh_wire_1834[ 30 ];
	assign fresh_wire_1888[ 31 ] = fresh_wire_1834[ 31 ];
	assign fresh_wire_1888[ 32 ] = fresh_wire_1834[ 32 ];
	assign fresh_wire_1888[ 33 ] = fresh_wire_1834[ 33 ];
	assign fresh_wire_1888[ 34 ] = fresh_wire_1834[ 34 ];
	assign fresh_wire_1888[ 35 ] = fresh_wire_1834[ 35 ];
	assign fresh_wire_1888[ 36 ] = fresh_wire_1834[ 36 ];
	assign fresh_wire_1888[ 37 ] = fresh_wire_1834[ 37 ];
	assign fresh_wire_1888[ 38 ] = fresh_wire_1834[ 38 ];
	assign fresh_wire_1888[ 39 ] = fresh_wire_1834[ 39 ];
	assign fresh_wire_1888[ 40 ] = fresh_wire_1834[ 40 ];
	assign fresh_wire_1888[ 41 ] = fresh_wire_1834[ 41 ];
	assign fresh_wire_1888[ 42 ] = fresh_wire_1834[ 42 ];
	assign fresh_wire_1888[ 43 ] = fresh_wire_1834[ 43 ];
	assign fresh_wire_1888[ 44 ] = fresh_wire_1834[ 44 ];
	assign fresh_wire_1888[ 45 ] = fresh_wire_1834[ 45 ];
	assign fresh_wire_1888[ 46 ] = fresh_wire_1834[ 46 ];
	assign fresh_wire_1888[ 47 ] = fresh_wire_1834[ 47 ];
	assign fresh_wire_1889[ 0 ] = fresh_wire_1572[ 0 ];
	assign fresh_wire_1889[ 1 ] = fresh_wire_1572[ 1 ];
	assign fresh_wire_1889[ 2 ] = fresh_wire_1572[ 2 ];
	assign fresh_wire_1889[ 3 ] = fresh_wire_1572[ 3 ];
	assign fresh_wire_1889[ 4 ] = fresh_wire_1572[ 4 ];
	assign fresh_wire_1889[ 5 ] = fresh_wire_1572[ 5 ];
	assign fresh_wire_1889[ 6 ] = fresh_wire_1572[ 6 ];
	assign fresh_wire_1889[ 7 ] = fresh_wire_1572[ 7 ];
	assign fresh_wire_1889[ 8 ] = fresh_wire_1572[ 8 ];
	assign fresh_wire_1889[ 9 ] = fresh_wire_1572[ 9 ];
	assign fresh_wire_1889[ 10 ] = fresh_wire_1572[ 10 ];
	assign fresh_wire_1889[ 11 ] = fresh_wire_1572[ 11 ];
	assign fresh_wire_1889[ 12 ] = fresh_wire_1572[ 12 ];
	assign fresh_wire_1889[ 13 ] = fresh_wire_1572[ 13 ];
	assign fresh_wire_1889[ 14 ] = fresh_wire_1572[ 14 ];
	assign fresh_wire_1889[ 15 ] = fresh_wire_1572[ 15 ];
	assign fresh_wire_1889[ 16 ] = fresh_wire_1834[ 0 ];
	assign fresh_wire_1889[ 17 ] = fresh_wire_1834[ 1 ];
	assign fresh_wire_1889[ 18 ] = fresh_wire_1834[ 2 ];
	assign fresh_wire_1889[ 19 ] = fresh_wire_1834[ 3 ];
	assign fresh_wire_1889[ 20 ] = fresh_wire_1834[ 4 ];
	assign fresh_wire_1889[ 21 ] = fresh_wire_1834[ 5 ];
	assign fresh_wire_1889[ 22 ] = fresh_wire_1834[ 6 ];
	assign fresh_wire_1889[ 23 ] = fresh_wire_1834[ 7 ];
	assign fresh_wire_1889[ 24 ] = fresh_wire_1834[ 8 ];
	assign fresh_wire_1889[ 25 ] = fresh_wire_1834[ 9 ];
	assign fresh_wire_1889[ 26 ] = fresh_wire_1834[ 10 ];
	assign fresh_wire_1889[ 27 ] = fresh_wire_1834[ 11 ];
	assign fresh_wire_1889[ 28 ] = fresh_wire_1834[ 12 ];
	assign fresh_wire_1889[ 29 ] = fresh_wire_1834[ 13 ];
	assign fresh_wire_1889[ 30 ] = fresh_wire_1834[ 14 ];
	assign fresh_wire_1889[ 31 ] = fresh_wire_1834[ 15 ];
	assign fresh_wire_1889[ 32 ] = fresh_wire_1834[ 16 ];
	assign fresh_wire_1889[ 33 ] = fresh_wire_1834[ 17 ];
	assign fresh_wire_1889[ 34 ] = fresh_wire_1834[ 18 ];
	assign fresh_wire_1889[ 35 ] = fresh_wire_1834[ 19 ];
	assign fresh_wire_1889[ 36 ] = fresh_wire_1834[ 20 ];
	assign fresh_wire_1889[ 37 ] = fresh_wire_1834[ 21 ];
	assign fresh_wire_1889[ 38 ] = fresh_wire_1834[ 22 ];
	assign fresh_wire_1889[ 39 ] = fresh_wire_1834[ 23 ];
	assign fresh_wire_1889[ 40 ] = fresh_wire_1834[ 24 ];
	assign fresh_wire_1889[ 41 ] = fresh_wire_1834[ 25 ];
	assign fresh_wire_1889[ 42 ] = fresh_wire_1834[ 26 ];
	assign fresh_wire_1889[ 43 ] = fresh_wire_1834[ 27 ];
	assign fresh_wire_1889[ 44 ] = fresh_wire_1834[ 28 ];
	assign fresh_wire_1889[ 45 ] = fresh_wire_1834[ 29 ];
	assign fresh_wire_1889[ 46 ] = fresh_wire_1834[ 30 ];
	assign fresh_wire_1889[ 47 ] = fresh_wire_1834[ 31 ];
	assign fresh_wire_1891[ 0 ] = fresh_wire_1700[ 0 ];
	assign fresh_wire_1892[ 0 ] = fresh_wire_1890[ 0 ];
	assign fresh_wire_1892[ 1 ] = fresh_wire_1890[ 1 ];
	assign fresh_wire_1892[ 2 ] = fresh_wire_1890[ 2 ];
	assign fresh_wire_1892[ 3 ] = fresh_wire_1890[ 3 ];
	assign fresh_wire_1892[ 4 ] = fresh_wire_1890[ 4 ];
	assign fresh_wire_1892[ 5 ] = fresh_wire_1890[ 5 ];
	assign fresh_wire_1892[ 6 ] = fresh_wire_1890[ 6 ];
	assign fresh_wire_1892[ 7 ] = fresh_wire_1890[ 7 ];
	assign fresh_wire_1892[ 8 ] = fresh_wire_1890[ 8 ];
	assign fresh_wire_1892[ 9 ] = fresh_wire_1890[ 9 ];
	assign fresh_wire_1892[ 10 ] = fresh_wire_1890[ 10 ];
	assign fresh_wire_1892[ 11 ] = fresh_wire_1890[ 11 ];
	assign fresh_wire_1892[ 12 ] = fresh_wire_1890[ 12 ];
	assign fresh_wire_1892[ 13 ] = fresh_wire_1890[ 13 ];
	assign fresh_wire_1892[ 14 ] = fresh_wire_1890[ 14 ];
	assign fresh_wire_1892[ 15 ] = fresh_wire_1890[ 15 ];
	assign fresh_wire_1892[ 16 ] = fresh_wire_1890[ 16 ];
	assign fresh_wire_1892[ 17 ] = fresh_wire_1890[ 17 ];
	assign fresh_wire_1892[ 18 ] = fresh_wire_1890[ 18 ];
	assign fresh_wire_1892[ 19 ] = fresh_wire_1890[ 19 ];
	assign fresh_wire_1892[ 20 ] = fresh_wire_1890[ 20 ];
	assign fresh_wire_1892[ 21 ] = fresh_wire_1890[ 21 ];
	assign fresh_wire_1892[ 22 ] = fresh_wire_1890[ 22 ];
	assign fresh_wire_1892[ 23 ] = fresh_wire_1890[ 23 ];
	assign fresh_wire_1892[ 24 ] = fresh_wire_1890[ 24 ];
	assign fresh_wire_1892[ 25 ] = fresh_wire_1890[ 25 ];
	assign fresh_wire_1892[ 26 ] = fresh_wire_1890[ 26 ];
	assign fresh_wire_1892[ 27 ] = fresh_wire_1890[ 27 ];
	assign fresh_wire_1892[ 28 ] = fresh_wire_1890[ 28 ];
	assign fresh_wire_1892[ 29 ] = fresh_wire_1890[ 29 ];
	assign fresh_wire_1892[ 30 ] = fresh_wire_1890[ 30 ];
	assign fresh_wire_1892[ 31 ] = fresh_wire_1890[ 31 ];
	assign fresh_wire_1892[ 32 ] = fresh_wire_1890[ 32 ];
	assign fresh_wire_1892[ 33 ] = fresh_wire_1890[ 33 ];
	assign fresh_wire_1892[ 34 ] = fresh_wire_1890[ 34 ];
	assign fresh_wire_1892[ 35 ] = fresh_wire_1890[ 35 ];
	assign fresh_wire_1892[ 36 ] = fresh_wire_1890[ 36 ];
	assign fresh_wire_1892[ 37 ] = fresh_wire_1890[ 37 ];
	assign fresh_wire_1892[ 38 ] = fresh_wire_1890[ 38 ];
	assign fresh_wire_1892[ 39 ] = fresh_wire_1890[ 39 ];
	assign fresh_wire_1892[ 40 ] = fresh_wire_1890[ 40 ];
	assign fresh_wire_1892[ 41 ] = fresh_wire_1890[ 41 ];
	assign fresh_wire_1892[ 42 ] = fresh_wire_1890[ 42 ];
	assign fresh_wire_1892[ 43 ] = fresh_wire_1890[ 43 ];
	assign fresh_wire_1892[ 44 ] = fresh_wire_1890[ 44 ];
	assign fresh_wire_1892[ 45 ] = fresh_wire_1890[ 45 ];
	assign fresh_wire_1892[ 46 ] = fresh_wire_1890[ 46 ];
	assign fresh_wire_1892[ 47 ] = fresh_wire_1890[ 47 ];
	assign fresh_wire_1893[ 0 ] = fresh_wire_1572[ 0 ];
	assign fresh_wire_1893[ 1 ] = fresh_wire_1572[ 1 ];
	assign fresh_wire_1893[ 2 ] = fresh_wire_1572[ 2 ];
	assign fresh_wire_1893[ 3 ] = fresh_wire_1572[ 3 ];
	assign fresh_wire_1893[ 4 ] = fresh_wire_1572[ 4 ];
	assign fresh_wire_1893[ 5 ] = fresh_wire_1572[ 5 ];
	assign fresh_wire_1893[ 6 ] = fresh_wire_1572[ 6 ];
	assign fresh_wire_1893[ 7 ] = fresh_wire_1572[ 7 ];
	assign fresh_wire_1893[ 8 ] = fresh_wire_1572[ 8 ];
	assign fresh_wire_1893[ 9 ] = fresh_wire_1572[ 9 ];
	assign fresh_wire_1893[ 10 ] = fresh_wire_1572[ 10 ];
	assign fresh_wire_1893[ 11 ] = fresh_wire_1572[ 11 ];
	assign fresh_wire_1893[ 12 ] = fresh_wire_1572[ 12 ];
	assign fresh_wire_1893[ 13 ] = fresh_wire_1572[ 13 ];
	assign fresh_wire_1893[ 14 ] = fresh_wire_1572[ 14 ];
	assign fresh_wire_1893[ 15 ] = fresh_wire_1572[ 15 ];
	assign fresh_wire_1893[ 16 ] = fresh_wire_1572[ 16 ];
	assign fresh_wire_1893[ 17 ] = fresh_wire_1572[ 17 ];
	assign fresh_wire_1893[ 18 ] = fresh_wire_1572[ 18 ];
	assign fresh_wire_1893[ 19 ] = fresh_wire_1572[ 19 ];
	assign fresh_wire_1893[ 20 ] = fresh_wire_1572[ 20 ];
	assign fresh_wire_1893[ 21 ] = fresh_wire_1572[ 21 ];
	assign fresh_wire_1893[ 22 ] = fresh_wire_1572[ 22 ];
	assign fresh_wire_1893[ 23 ] = fresh_wire_1572[ 23 ];
	assign fresh_wire_1893[ 24 ] = fresh_wire_1572[ 24 ];
	assign fresh_wire_1893[ 25 ] = fresh_wire_1572[ 25 ];
	assign fresh_wire_1893[ 26 ] = fresh_wire_1572[ 26 ];
	assign fresh_wire_1893[ 27 ] = fresh_wire_1572[ 27 ];
	assign fresh_wire_1893[ 28 ] = fresh_wire_1572[ 28 ];
	assign fresh_wire_1893[ 29 ] = fresh_wire_1572[ 29 ];
	assign fresh_wire_1893[ 30 ] = fresh_wire_1572[ 30 ];
	assign fresh_wire_1893[ 31 ] = fresh_wire_1572[ 31 ];
	assign fresh_wire_1893[ 32 ] = fresh_wire_1834[ 0 ];
	assign fresh_wire_1893[ 33 ] = fresh_wire_1834[ 1 ];
	assign fresh_wire_1893[ 34 ] = fresh_wire_1834[ 2 ];
	assign fresh_wire_1893[ 35 ] = fresh_wire_1834[ 3 ];
	assign fresh_wire_1893[ 36 ] = fresh_wire_1834[ 4 ];
	assign fresh_wire_1893[ 37 ] = fresh_wire_1834[ 5 ];
	assign fresh_wire_1893[ 38 ] = fresh_wire_1834[ 6 ];
	assign fresh_wire_1893[ 39 ] = fresh_wire_1834[ 7 ];
	assign fresh_wire_1893[ 40 ] = fresh_wire_1834[ 8 ];
	assign fresh_wire_1893[ 41 ] = fresh_wire_1834[ 9 ];
	assign fresh_wire_1893[ 42 ] = fresh_wire_1834[ 10 ];
	assign fresh_wire_1893[ 43 ] = fresh_wire_1834[ 11 ];
	assign fresh_wire_1893[ 44 ] = fresh_wire_1834[ 12 ];
	assign fresh_wire_1893[ 45 ] = fresh_wire_1834[ 13 ];
	assign fresh_wire_1893[ 46 ] = fresh_wire_1834[ 14 ];
	assign fresh_wire_1893[ 47 ] = fresh_wire_1834[ 15 ];
	assign fresh_wire_1895[ 0 ] = fresh_wire_1706[ 0 ];
	assign fresh_wire_1896[ 0 ] = fresh_wire_1830[ 0 ];
	assign fresh_wire_1896[ 1 ] = fresh_wire_1830[ 1 ];
	assign fresh_wire_1897[ 0 ] = fresh_wire_1899[ 0 ];
	assign fresh_wire_1897[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1900[ 0 ] = fresh_wire_1129[ 0 ];
	assign fresh_wire_1902[ 0 ] = fresh_wire_1398[ 0 ];
	assign fresh_wire_1904[ 0 ] = fresh_wire_1901[ 0 ];
	assign fresh_wire_1905[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1907[ 0 ] = fresh_wire_1903[ 0 ];
	assign fresh_wire_1908[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1910[ 0 ] = fresh_wire_1915[ 0 ];
	assign fresh_wire_1910[ 1 ] = fresh_wire_1915[ 1 ];
	assign fresh_wire_1910[ 2 ] = fresh_wire_1915[ 2 ];
	assign fresh_wire_1910[ 3 ] = fresh_wire_1915[ 3 ];
	assign fresh_wire_1910[ 4 ] = fresh_wire_1915[ 4 ];
	assign fresh_wire_1910[ 5 ] = fresh_wire_1915[ 5 ];
	assign fresh_wire_1910[ 6 ] = fresh_wire_1915[ 6 ];
	assign fresh_wire_1910[ 7 ] = fresh_wire_1915[ 7 ];
	assign fresh_wire_1910[ 8 ] = fresh_wire_1915[ 8 ];
	assign fresh_wire_1910[ 9 ] = fresh_wire_1915[ 9 ];
	assign fresh_wire_1910[ 10 ] = fresh_wire_1915[ 10 ];
	assign fresh_wire_1910[ 11 ] = fresh_wire_1915[ 11 ];
	assign fresh_wire_1910[ 12 ] = fresh_wire_1915[ 12 ];
	assign fresh_wire_1910[ 13 ] = fresh_wire_1915[ 13 ];
	assign fresh_wire_1910[ 14 ] = fresh_wire_1915[ 14 ];
	assign fresh_wire_1910[ 15 ] = fresh_wire_1915[ 15 ];
	assign fresh_wire_1912[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1913[ 0 ] = fresh_wire_1911[ 0 ];
	assign fresh_wire_1913[ 1 ] = fresh_wire_1911[ 1 ];
	assign fresh_wire_1913[ 2 ] = fresh_wire_1911[ 2 ];
	assign fresh_wire_1913[ 3 ] = fresh_wire_1911[ 3 ];
	assign fresh_wire_1913[ 4 ] = fresh_wire_1911[ 4 ];
	assign fresh_wire_1913[ 5 ] = fresh_wire_1911[ 5 ];
	assign fresh_wire_1913[ 6 ] = fresh_wire_1911[ 6 ];
	assign fresh_wire_1913[ 7 ] = fresh_wire_1911[ 7 ];
	assign fresh_wire_1913[ 8 ] = fresh_wire_1911[ 8 ];
	assign fresh_wire_1913[ 9 ] = fresh_wire_1911[ 9 ];
	assign fresh_wire_1913[ 10 ] = fresh_wire_1911[ 10 ];
	assign fresh_wire_1913[ 11 ] = fresh_wire_1911[ 11 ];
	assign fresh_wire_1913[ 12 ] = fresh_wire_1911[ 12 ];
	assign fresh_wire_1913[ 13 ] = fresh_wire_1911[ 13 ];
	assign fresh_wire_1913[ 14 ] = fresh_wire_1911[ 14 ];
	assign fresh_wire_1913[ 15 ] = fresh_wire_1911[ 15 ];
	assign fresh_wire_1914[ 0 ] = fresh_wire_1994[ 0 ];
	assign fresh_wire_1914[ 1 ] = fresh_wire_1994[ 1 ];
	assign fresh_wire_1914[ 2 ] = fresh_wire_1994[ 2 ];
	assign fresh_wire_1914[ 3 ] = fresh_wire_1994[ 3 ];
	assign fresh_wire_1914[ 4 ] = fresh_wire_1994[ 4 ];
	assign fresh_wire_1914[ 5 ] = fresh_wire_1994[ 5 ];
	assign fresh_wire_1914[ 6 ] = fresh_wire_1994[ 6 ];
	assign fresh_wire_1914[ 7 ] = fresh_wire_1994[ 7 ];
	assign fresh_wire_1914[ 8 ] = fresh_wire_1994[ 8 ];
	assign fresh_wire_1914[ 9 ] = fresh_wire_1994[ 9 ];
	assign fresh_wire_1914[ 10 ] = fresh_wire_1994[ 10 ];
	assign fresh_wire_1914[ 11 ] = fresh_wire_1994[ 11 ];
	assign fresh_wire_1914[ 12 ] = fresh_wire_1994[ 12 ];
	assign fresh_wire_1914[ 13 ] = fresh_wire_1994[ 13 ];
	assign fresh_wire_1914[ 14 ] = fresh_wire_1994[ 14 ];
	assign fresh_wire_1914[ 15 ] = fresh_wire_1994[ 15 ];
	assign fresh_wire_1916[ 0 ] = fresh_wire_1906[ 0 ];
	assign fresh_wire_1917[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1917[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1917[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1917[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1917[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1917[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1917[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1917[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1917[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1917[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1917[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1917[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1917[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1917[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1917[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1917[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1918[ 0 ] = fresh_wire_1921[ 0 ];
	assign fresh_wire_1918[ 1 ] = fresh_wire_1921[ 0 ];
	assign fresh_wire_1918[ 2 ] = fresh_wire_1921[ 0 ];
	assign fresh_wire_1918[ 3 ] = fresh_wire_1921[ 0 ];
	assign fresh_wire_1918[ 4 ] = fresh_wire_1921[ 0 ];
	assign fresh_wire_1918[ 5 ] = fresh_wire_1921[ 0 ];
	assign fresh_wire_1918[ 6 ] = fresh_wire_1921[ 0 ];
	assign fresh_wire_1918[ 7 ] = fresh_wire_1921[ 0 ];
	assign fresh_wire_1918[ 8 ] = fresh_wire_1921[ 0 ];
	assign fresh_wire_1918[ 9 ] = fresh_wire_1921[ 0 ];
	assign fresh_wire_1918[ 10 ] = fresh_wire_1921[ 0 ];
	assign fresh_wire_1918[ 11 ] = fresh_wire_1921[ 0 ];
	assign fresh_wire_1918[ 12 ] = fresh_wire_1921[ 0 ];
	assign fresh_wire_1918[ 13 ] = fresh_wire_1921[ 0 ];
	assign fresh_wire_1918[ 14 ] = fresh_wire_1921[ 0 ];
	assign fresh_wire_1918[ 15 ] = fresh_wire_1921[ 0 ];
	assign fresh_wire_1920[ 0 ] = fresh_wire_1909[ 0 ];
	assign fresh_wire_1922[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1922[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1922[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1922[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1922[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1922[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1922[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1922[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1922[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1922[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1922[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1922[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1922[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1922[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1922[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1922[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_1923[ 0 ] = fresh_wire_1919[ 0 ];
	assign fresh_wire_1923[ 1 ] = fresh_wire_1919[ 1 ];
	assign fresh_wire_1923[ 2 ] = fresh_wire_1919[ 2 ];
	assign fresh_wire_1923[ 3 ] = fresh_wire_1919[ 3 ];
	assign fresh_wire_1923[ 4 ] = fresh_wire_1919[ 4 ];
	assign fresh_wire_1923[ 5 ] = fresh_wire_1919[ 5 ];
	assign fresh_wire_1923[ 6 ] = fresh_wire_1919[ 6 ];
	assign fresh_wire_1923[ 7 ] = fresh_wire_1919[ 7 ];
	assign fresh_wire_1923[ 8 ] = fresh_wire_1919[ 8 ];
	assign fresh_wire_1923[ 9 ] = fresh_wire_1919[ 9 ];
	assign fresh_wire_1923[ 10 ] = fresh_wire_1919[ 10 ];
	assign fresh_wire_1923[ 11 ] = fresh_wire_1919[ 11 ];
	assign fresh_wire_1923[ 12 ] = fresh_wire_1919[ 12 ];
	assign fresh_wire_1923[ 13 ] = fresh_wire_1919[ 13 ];
	assign fresh_wire_1923[ 14 ] = fresh_wire_1919[ 14 ];
	assign fresh_wire_1923[ 15 ] = fresh_wire_1919[ 15 ];
	assign fresh_wire_1925[ 0 ] = fresh_wire_1906[ 0 ];
	assign fresh_wire_1926[ 0 ] = fresh_wire_1930[ 0 ];
	assign fresh_wire_1926[ 1 ] = fresh_wire_1937[ 0 ];
	assign fresh_wire_1926[ 2 ] = fresh_wire_1938[ 0 ];
	assign fresh_wire_1926[ 3 ] = fresh_wire_1939[ 0 ];
	assign fresh_wire_1926[ 4 ] = fresh_wire_1940[ 0 ];
	assign fresh_wire_1926[ 5 ] = fresh_wire_1941[ 0 ];
	assign fresh_wire_1926[ 6 ] = fresh_wire_1942[ 0 ];
	assign fresh_wire_1926[ 7 ] = fresh_wire_1943[ 0 ];
	assign fresh_wire_1926[ 8 ] = fresh_wire_1944[ 0 ];
	assign fresh_wire_1926[ 9 ] = fresh_wire_1945[ 0 ];
	assign fresh_wire_1926[ 10 ] = fresh_wire_1931[ 0 ];
	assign fresh_wire_1926[ 11 ] = fresh_wire_1932[ 0 ];
	assign fresh_wire_1926[ 12 ] = fresh_wire_1933[ 0 ];
	assign fresh_wire_1926[ 13 ] = fresh_wire_1934[ 0 ];
	assign fresh_wire_1926[ 14 ] = fresh_wire_1935[ 0 ];
	assign fresh_wire_1926[ 15 ] = fresh_wire_1936[ 0 ];
	assign fresh_wire_1927[ 0 ] = fresh_wire_1686[ 0 ];
	assign fresh_wire_1927[ 1 ] = fresh_wire_1686[ 1 ];
	assign fresh_wire_1927[ 2 ] = fresh_wire_1686[ 2 ];
	assign fresh_wire_1927[ 3 ] = fresh_wire_1686[ 3 ];
	assign fresh_wire_1927[ 4 ] = fresh_wire_1686[ 4 ];
	assign fresh_wire_1927[ 5 ] = fresh_wire_1686[ 5 ];
	assign fresh_wire_1927[ 6 ] = fresh_wire_1686[ 6 ];
	assign fresh_wire_1927[ 7 ] = fresh_wire_1686[ 7 ];
	assign fresh_wire_1927[ 8 ] = fresh_wire_1686[ 8 ];
	assign fresh_wire_1927[ 9 ] = fresh_wire_1686[ 9 ];
	assign fresh_wire_1927[ 10 ] = fresh_wire_1686[ 10 ];
	assign fresh_wire_1927[ 11 ] = fresh_wire_1686[ 11 ];
	assign fresh_wire_1927[ 12 ] = fresh_wire_1686[ 12 ];
	assign fresh_wire_1927[ 13 ] = fresh_wire_1686[ 13 ];
	assign fresh_wire_1927[ 14 ] = fresh_wire_1686[ 14 ];
	assign fresh_wire_1927[ 15 ] = fresh_wire_1686[ 15 ];
	assign fresh_wire_1929[ 0 ] = fresh_wire_1909[ 0 ];
	assign fresh_wire_1946[ 0 ] = fresh_wire_1950[ 0 ];
	assign fresh_wire_1946[ 1 ] = fresh_wire_1957[ 0 ];
	assign fresh_wire_1946[ 2 ] = fresh_wire_1958[ 0 ];
	assign fresh_wire_1946[ 3 ] = fresh_wire_1959[ 0 ];
	assign fresh_wire_1946[ 4 ] = fresh_wire_1960[ 0 ];
	assign fresh_wire_1946[ 5 ] = fresh_wire_1961[ 0 ];
	assign fresh_wire_1946[ 6 ] = fresh_wire_1962[ 0 ];
	assign fresh_wire_1946[ 7 ] = fresh_wire_1963[ 0 ];
	assign fresh_wire_1946[ 8 ] = fresh_wire_1964[ 0 ];
	assign fresh_wire_1946[ 9 ] = fresh_wire_1965[ 0 ];
	assign fresh_wire_1946[ 10 ] = fresh_wire_1951[ 0 ];
	assign fresh_wire_1946[ 11 ] = fresh_wire_1952[ 0 ];
	assign fresh_wire_1946[ 12 ] = fresh_wire_1953[ 0 ];
	assign fresh_wire_1946[ 13 ] = fresh_wire_1954[ 0 ];
	assign fresh_wire_1946[ 14 ] = fresh_wire_1955[ 0 ];
	assign fresh_wire_1946[ 15 ] = fresh_wire_1956[ 0 ];
	assign fresh_wire_1947[ 0 ] = fresh_wire_1928[ 0 ];
	assign fresh_wire_1947[ 1 ] = fresh_wire_1928[ 1 ];
	assign fresh_wire_1947[ 2 ] = fresh_wire_1928[ 2 ];
	assign fresh_wire_1947[ 3 ] = fresh_wire_1928[ 3 ];
	assign fresh_wire_1947[ 4 ] = fresh_wire_1928[ 4 ];
	assign fresh_wire_1947[ 5 ] = fresh_wire_1928[ 5 ];
	assign fresh_wire_1947[ 6 ] = fresh_wire_1928[ 6 ];
	assign fresh_wire_1947[ 7 ] = fresh_wire_1928[ 7 ];
	assign fresh_wire_1947[ 8 ] = fresh_wire_1928[ 8 ];
	assign fresh_wire_1947[ 9 ] = fresh_wire_1928[ 9 ];
	assign fresh_wire_1947[ 10 ] = fresh_wire_1928[ 10 ];
	assign fresh_wire_1947[ 11 ] = fresh_wire_1928[ 11 ];
	assign fresh_wire_1947[ 12 ] = fresh_wire_1928[ 12 ];
	assign fresh_wire_1947[ 13 ] = fresh_wire_1928[ 13 ];
	assign fresh_wire_1947[ 14 ] = fresh_wire_1928[ 14 ];
	assign fresh_wire_1947[ 15 ] = fresh_wire_1928[ 15 ];
	assign fresh_wire_1949[ 0 ] = fresh_wire_1906[ 0 ];
	assign fresh_wire_1966[ 0 ] = fresh_wire_1970[ 0 ];
	assign fresh_wire_1966[ 1 ] = fresh_wire_1971[ 0 ];
	assign fresh_wire_1966[ 2 ] = fresh_wire_1972[ 0 ];
	assign fresh_wire_1966[ 3 ] = fresh_wire_1973[ 0 ];
	assign fresh_wire_1966[ 4 ] = fresh_wire_1974[ 0 ];
	assign fresh_wire_1966[ 5 ] = fresh_wire_1975[ 0 ];
	assign fresh_wire_1966[ 6 ] = fresh_wire_1976[ 0 ];
	assign fresh_wire_1966[ 7 ] = fresh_wire_1977[ 0 ];
	assign fresh_wire_1966[ 8 ] = fresh_wire_1978[ 0 ];
	assign fresh_wire_1967[ 0 ] = fresh_wire_1407[ 0 ];
	assign fresh_wire_1967[ 1 ] = fresh_wire_1407[ 1 ];
	assign fresh_wire_1967[ 2 ] = fresh_wire_1407[ 2 ];
	assign fresh_wire_1967[ 3 ] = fresh_wire_1407[ 3 ];
	assign fresh_wire_1967[ 4 ] = fresh_wire_1407[ 4 ];
	assign fresh_wire_1967[ 5 ] = fresh_wire_1407[ 5 ];
	assign fresh_wire_1967[ 6 ] = fresh_wire_1407[ 6 ];
	assign fresh_wire_1967[ 7 ] = fresh_wire_1407[ 7 ];
	assign fresh_wire_1967[ 8 ] = fresh_wire_1407[ 8 ];
	assign fresh_wire_1969[ 0 ] = fresh_wire_1909[ 0 ];
	assign fresh_wire_1979[ 0 ] = fresh_wire_1983[ 0 ];
	assign fresh_wire_1979[ 1 ] = fresh_wire_1984[ 0 ];
	assign fresh_wire_1979[ 2 ] = fresh_wire_1985[ 0 ];
	assign fresh_wire_1979[ 3 ] = fresh_wire_1986[ 0 ];
	assign fresh_wire_1979[ 4 ] = fresh_wire_1987[ 0 ];
	assign fresh_wire_1979[ 5 ] = fresh_wire_1988[ 0 ];
	assign fresh_wire_1979[ 6 ] = fresh_wire_1989[ 0 ];
	assign fresh_wire_1979[ 7 ] = fresh_wire_1990[ 0 ];
	assign fresh_wire_1979[ 8 ] = fresh_wire_1991[ 0 ];
	assign fresh_wire_1980[ 0 ] = fresh_wire_1968[ 0 ];
	assign fresh_wire_1980[ 1 ] = fresh_wire_1968[ 1 ];
	assign fresh_wire_1980[ 2 ] = fresh_wire_1968[ 2 ];
	assign fresh_wire_1980[ 3 ] = fresh_wire_1968[ 3 ];
	assign fresh_wire_1980[ 4 ] = fresh_wire_1968[ 4 ];
	assign fresh_wire_1980[ 5 ] = fresh_wire_1968[ 5 ];
	assign fresh_wire_1980[ 6 ] = fresh_wire_1968[ 6 ];
	assign fresh_wire_1980[ 7 ] = fresh_wire_1968[ 7 ];
	assign fresh_wire_1980[ 8 ] = fresh_wire_1968[ 8 ];
	assign fresh_wire_1982[ 0 ] = fresh_wire_1906[ 0 ];
	assign fresh_wire_1992[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_1993[ 0 ] = fresh_wire_1407[ 0 ];
	assign fresh_wire_1993[ 1 ] = fresh_wire_1407[ 1 ];
	assign fresh_wire_1993[ 2 ] = fresh_wire_1407[ 2 ];
	assign fresh_wire_1993[ 3 ] = fresh_wire_1407[ 3 ];
	assign fresh_wire_1993[ 4 ] = fresh_wire_1407[ 4 ];
	assign fresh_wire_1993[ 5 ] = fresh_wire_1407[ 5 ];
	assign fresh_wire_1993[ 6 ] = fresh_wire_1407[ 6 ];
	assign fresh_wire_1993[ 7 ] = fresh_wire_1407[ 7 ];
	assign fresh_wire_1993[ 8 ] = fresh_wire_1407[ 8 ];
	assign fresh_wire_1995[ 0 ] = fresh_wire_1981[ 0 ];
	assign fresh_wire_1995[ 1 ] = fresh_wire_1981[ 1 ];
	assign fresh_wire_1995[ 2 ] = fresh_wire_1981[ 2 ];
	assign fresh_wire_1995[ 3 ] = fresh_wire_1981[ 3 ];
	assign fresh_wire_1995[ 4 ] = fresh_wire_1981[ 4 ];
	assign fresh_wire_1995[ 5 ] = fresh_wire_1981[ 5 ];
	assign fresh_wire_1995[ 6 ] = fresh_wire_1981[ 6 ];
	assign fresh_wire_1995[ 7 ] = fresh_wire_1981[ 7 ];
	assign fresh_wire_1995[ 8 ] = fresh_wire_1981[ 8 ];
	assign fresh_wire_1996[ 0 ] = fresh_wire_1948[ 0 ];
	assign fresh_wire_1996[ 1 ] = fresh_wire_1948[ 1 ];
	assign fresh_wire_1996[ 2 ] = fresh_wire_1948[ 2 ];
	assign fresh_wire_1996[ 3 ] = fresh_wire_1948[ 3 ];
	assign fresh_wire_1996[ 4 ] = fresh_wire_1948[ 4 ];
	assign fresh_wire_1996[ 5 ] = fresh_wire_1948[ 5 ];
	assign fresh_wire_1996[ 6 ] = fresh_wire_1948[ 6 ];
	assign fresh_wire_1996[ 7 ] = fresh_wire_1948[ 7 ];
	assign fresh_wire_1996[ 8 ] = fresh_wire_1948[ 8 ];
	assign fresh_wire_1996[ 9 ] = fresh_wire_1948[ 9 ];
	assign fresh_wire_1996[ 10 ] = fresh_wire_1948[ 10 ];
	assign fresh_wire_1996[ 11 ] = fresh_wire_1948[ 11 ];
	assign fresh_wire_1996[ 12 ] = fresh_wire_1948[ 12 ];
	assign fresh_wire_1996[ 13 ] = fresh_wire_1948[ 13 ];
	assign fresh_wire_1996[ 14 ] = fresh_wire_1948[ 14 ];
	assign fresh_wire_1996[ 15 ] = fresh_wire_1948[ 15 ];
	assign fresh_wire_1997[ 0 ] = fresh_wire_1924[ 0 ];
	assign fresh_wire_1998[ 0 ] = fresh_wire_1132[ 0 ];
	assign fresh_wire_2000[ 0 ] = fresh_wire_1398[ 0 ];
	assign fresh_wire_2002[ 0 ] = fresh_wire_1999[ 0 ];
	assign fresh_wire_2003[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2005[ 0 ] = fresh_wire_2001[ 0 ];
	assign fresh_wire_2006[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2008[ 0 ] = fresh_wire_2013[ 0 ];
	assign fresh_wire_2008[ 1 ] = fresh_wire_2013[ 1 ];
	assign fresh_wire_2008[ 2 ] = fresh_wire_2013[ 2 ];
	assign fresh_wire_2008[ 3 ] = fresh_wire_2013[ 3 ];
	assign fresh_wire_2008[ 4 ] = fresh_wire_2013[ 4 ];
	assign fresh_wire_2008[ 5 ] = fresh_wire_2013[ 5 ];
	assign fresh_wire_2008[ 6 ] = fresh_wire_2013[ 6 ];
	assign fresh_wire_2008[ 7 ] = fresh_wire_2013[ 7 ];
	assign fresh_wire_2008[ 8 ] = fresh_wire_2013[ 8 ];
	assign fresh_wire_2008[ 9 ] = fresh_wire_2013[ 9 ];
	assign fresh_wire_2008[ 10 ] = fresh_wire_2013[ 10 ];
	assign fresh_wire_2008[ 11 ] = fresh_wire_2013[ 11 ];
	assign fresh_wire_2008[ 12 ] = fresh_wire_2013[ 12 ];
	assign fresh_wire_2008[ 13 ] = fresh_wire_2013[ 13 ];
	assign fresh_wire_2008[ 14 ] = fresh_wire_2013[ 14 ];
	assign fresh_wire_2008[ 15 ] = fresh_wire_2013[ 15 ];
	assign fresh_wire_2010[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_2011[ 0 ] = fresh_wire_2009[ 0 ];
	assign fresh_wire_2011[ 1 ] = fresh_wire_2009[ 1 ];
	assign fresh_wire_2011[ 2 ] = fresh_wire_2009[ 2 ];
	assign fresh_wire_2011[ 3 ] = fresh_wire_2009[ 3 ];
	assign fresh_wire_2011[ 4 ] = fresh_wire_2009[ 4 ];
	assign fresh_wire_2011[ 5 ] = fresh_wire_2009[ 5 ];
	assign fresh_wire_2011[ 6 ] = fresh_wire_2009[ 6 ];
	assign fresh_wire_2011[ 7 ] = fresh_wire_2009[ 7 ];
	assign fresh_wire_2011[ 8 ] = fresh_wire_2009[ 8 ];
	assign fresh_wire_2011[ 9 ] = fresh_wire_2009[ 9 ];
	assign fresh_wire_2011[ 10 ] = fresh_wire_2009[ 10 ];
	assign fresh_wire_2011[ 11 ] = fresh_wire_2009[ 11 ];
	assign fresh_wire_2011[ 12 ] = fresh_wire_2009[ 12 ];
	assign fresh_wire_2011[ 13 ] = fresh_wire_2009[ 13 ];
	assign fresh_wire_2011[ 14 ] = fresh_wire_2009[ 14 ];
	assign fresh_wire_2011[ 15 ] = fresh_wire_2009[ 15 ];
	assign fresh_wire_2012[ 0 ] = fresh_wire_2092[ 0 ];
	assign fresh_wire_2012[ 1 ] = fresh_wire_2092[ 1 ];
	assign fresh_wire_2012[ 2 ] = fresh_wire_2092[ 2 ];
	assign fresh_wire_2012[ 3 ] = fresh_wire_2092[ 3 ];
	assign fresh_wire_2012[ 4 ] = fresh_wire_2092[ 4 ];
	assign fresh_wire_2012[ 5 ] = fresh_wire_2092[ 5 ];
	assign fresh_wire_2012[ 6 ] = fresh_wire_2092[ 6 ];
	assign fresh_wire_2012[ 7 ] = fresh_wire_2092[ 7 ];
	assign fresh_wire_2012[ 8 ] = fresh_wire_2092[ 8 ];
	assign fresh_wire_2012[ 9 ] = fresh_wire_2092[ 9 ];
	assign fresh_wire_2012[ 10 ] = fresh_wire_2092[ 10 ];
	assign fresh_wire_2012[ 11 ] = fresh_wire_2092[ 11 ];
	assign fresh_wire_2012[ 12 ] = fresh_wire_2092[ 12 ];
	assign fresh_wire_2012[ 13 ] = fresh_wire_2092[ 13 ];
	assign fresh_wire_2012[ 14 ] = fresh_wire_2092[ 14 ];
	assign fresh_wire_2012[ 15 ] = fresh_wire_2092[ 15 ];
	assign fresh_wire_2014[ 0 ] = fresh_wire_2004[ 0 ];
	assign fresh_wire_2015[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2015[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2015[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2015[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2015[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2015[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2015[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2015[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2015[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2015[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2015[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2015[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2015[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2015[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2015[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2015[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2016[ 0 ] = fresh_wire_2019[ 0 ];
	assign fresh_wire_2016[ 1 ] = fresh_wire_2019[ 0 ];
	assign fresh_wire_2016[ 2 ] = fresh_wire_2019[ 0 ];
	assign fresh_wire_2016[ 3 ] = fresh_wire_2019[ 0 ];
	assign fresh_wire_2016[ 4 ] = fresh_wire_2019[ 0 ];
	assign fresh_wire_2016[ 5 ] = fresh_wire_2019[ 0 ];
	assign fresh_wire_2016[ 6 ] = fresh_wire_2019[ 0 ];
	assign fresh_wire_2016[ 7 ] = fresh_wire_2019[ 0 ];
	assign fresh_wire_2016[ 8 ] = fresh_wire_2019[ 0 ];
	assign fresh_wire_2016[ 9 ] = fresh_wire_2019[ 0 ];
	assign fresh_wire_2016[ 10 ] = fresh_wire_2019[ 0 ];
	assign fresh_wire_2016[ 11 ] = fresh_wire_2019[ 0 ];
	assign fresh_wire_2016[ 12 ] = fresh_wire_2019[ 0 ];
	assign fresh_wire_2016[ 13 ] = fresh_wire_2019[ 0 ];
	assign fresh_wire_2016[ 14 ] = fresh_wire_2019[ 0 ];
	assign fresh_wire_2016[ 15 ] = fresh_wire_2019[ 0 ];
	assign fresh_wire_2018[ 0 ] = fresh_wire_2007[ 0 ];
	assign fresh_wire_2020[ 0 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2020[ 1 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2020[ 2 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2020[ 3 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2020[ 4 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2020[ 5 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2020[ 6 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2020[ 7 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2020[ 8 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2020[ 9 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2020[ 10 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2020[ 11 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2020[ 12 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2020[ 13 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2020[ 14 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2020[ 15 ] = fresh_wire_2249[ 0 ];
	assign fresh_wire_2021[ 0 ] = fresh_wire_2017[ 0 ];
	assign fresh_wire_2021[ 1 ] = fresh_wire_2017[ 1 ];
	assign fresh_wire_2021[ 2 ] = fresh_wire_2017[ 2 ];
	assign fresh_wire_2021[ 3 ] = fresh_wire_2017[ 3 ];
	assign fresh_wire_2021[ 4 ] = fresh_wire_2017[ 4 ];
	assign fresh_wire_2021[ 5 ] = fresh_wire_2017[ 5 ];
	assign fresh_wire_2021[ 6 ] = fresh_wire_2017[ 6 ];
	assign fresh_wire_2021[ 7 ] = fresh_wire_2017[ 7 ];
	assign fresh_wire_2021[ 8 ] = fresh_wire_2017[ 8 ];
	assign fresh_wire_2021[ 9 ] = fresh_wire_2017[ 9 ];
	assign fresh_wire_2021[ 10 ] = fresh_wire_2017[ 10 ];
	assign fresh_wire_2021[ 11 ] = fresh_wire_2017[ 11 ];
	assign fresh_wire_2021[ 12 ] = fresh_wire_2017[ 12 ];
	assign fresh_wire_2021[ 13 ] = fresh_wire_2017[ 13 ];
	assign fresh_wire_2021[ 14 ] = fresh_wire_2017[ 14 ];
	assign fresh_wire_2021[ 15 ] = fresh_wire_2017[ 15 ];
	assign fresh_wire_2023[ 0 ] = fresh_wire_2004[ 0 ];
	assign fresh_wire_2024[ 0 ] = fresh_wire_2028[ 0 ];
	assign fresh_wire_2024[ 1 ] = fresh_wire_2035[ 0 ];
	assign fresh_wire_2024[ 2 ] = fresh_wire_2036[ 0 ];
	assign fresh_wire_2024[ 3 ] = fresh_wire_2037[ 0 ];
	assign fresh_wire_2024[ 4 ] = fresh_wire_2038[ 0 ];
	assign fresh_wire_2024[ 5 ] = fresh_wire_2039[ 0 ];
	assign fresh_wire_2024[ 6 ] = fresh_wire_2040[ 0 ];
	assign fresh_wire_2024[ 7 ] = fresh_wire_2041[ 0 ];
	assign fresh_wire_2024[ 8 ] = fresh_wire_2042[ 0 ];
	assign fresh_wire_2024[ 9 ] = fresh_wire_2043[ 0 ];
	assign fresh_wire_2024[ 10 ] = fresh_wire_2029[ 0 ];
	assign fresh_wire_2024[ 11 ] = fresh_wire_2030[ 0 ];
	assign fresh_wire_2024[ 12 ] = fresh_wire_2031[ 0 ];
	assign fresh_wire_2024[ 13 ] = fresh_wire_2032[ 0 ];
	assign fresh_wire_2024[ 14 ] = fresh_wire_2033[ 0 ];
	assign fresh_wire_2024[ 15 ] = fresh_wire_2034[ 0 ];
	assign fresh_wire_2025[ 0 ] = fresh_wire_1686[ 16 ];
	assign fresh_wire_2025[ 1 ] = fresh_wire_1686[ 17 ];
	assign fresh_wire_2025[ 2 ] = fresh_wire_1686[ 18 ];
	assign fresh_wire_2025[ 3 ] = fresh_wire_1686[ 19 ];
	assign fresh_wire_2025[ 4 ] = fresh_wire_1686[ 20 ];
	assign fresh_wire_2025[ 5 ] = fresh_wire_1686[ 21 ];
	assign fresh_wire_2025[ 6 ] = fresh_wire_1686[ 22 ];
	assign fresh_wire_2025[ 7 ] = fresh_wire_1686[ 23 ];
	assign fresh_wire_2025[ 8 ] = fresh_wire_1686[ 24 ];
	assign fresh_wire_2025[ 9 ] = fresh_wire_1686[ 25 ];
	assign fresh_wire_2025[ 10 ] = fresh_wire_1686[ 26 ];
	assign fresh_wire_2025[ 11 ] = fresh_wire_1686[ 27 ];
	assign fresh_wire_2025[ 12 ] = fresh_wire_1686[ 28 ];
	assign fresh_wire_2025[ 13 ] = fresh_wire_1686[ 29 ];
	assign fresh_wire_2025[ 14 ] = fresh_wire_1686[ 30 ];
	assign fresh_wire_2025[ 15 ] = fresh_wire_1686[ 31 ];
	assign fresh_wire_2027[ 0 ] = fresh_wire_2007[ 0 ];
	assign fresh_wire_2044[ 0 ] = fresh_wire_2048[ 0 ];
	assign fresh_wire_2044[ 1 ] = fresh_wire_2055[ 0 ];
	assign fresh_wire_2044[ 2 ] = fresh_wire_2056[ 0 ];
	assign fresh_wire_2044[ 3 ] = fresh_wire_2057[ 0 ];
	assign fresh_wire_2044[ 4 ] = fresh_wire_2058[ 0 ];
	assign fresh_wire_2044[ 5 ] = fresh_wire_2059[ 0 ];
	assign fresh_wire_2044[ 6 ] = fresh_wire_2060[ 0 ];
	assign fresh_wire_2044[ 7 ] = fresh_wire_2061[ 0 ];
	assign fresh_wire_2044[ 8 ] = fresh_wire_2062[ 0 ];
	assign fresh_wire_2044[ 9 ] = fresh_wire_2063[ 0 ];
	assign fresh_wire_2044[ 10 ] = fresh_wire_2049[ 0 ];
	assign fresh_wire_2044[ 11 ] = fresh_wire_2050[ 0 ];
	assign fresh_wire_2044[ 12 ] = fresh_wire_2051[ 0 ];
	assign fresh_wire_2044[ 13 ] = fresh_wire_2052[ 0 ];
	assign fresh_wire_2044[ 14 ] = fresh_wire_2053[ 0 ];
	assign fresh_wire_2044[ 15 ] = fresh_wire_2054[ 0 ];
	assign fresh_wire_2045[ 0 ] = fresh_wire_2026[ 0 ];
	assign fresh_wire_2045[ 1 ] = fresh_wire_2026[ 1 ];
	assign fresh_wire_2045[ 2 ] = fresh_wire_2026[ 2 ];
	assign fresh_wire_2045[ 3 ] = fresh_wire_2026[ 3 ];
	assign fresh_wire_2045[ 4 ] = fresh_wire_2026[ 4 ];
	assign fresh_wire_2045[ 5 ] = fresh_wire_2026[ 5 ];
	assign fresh_wire_2045[ 6 ] = fresh_wire_2026[ 6 ];
	assign fresh_wire_2045[ 7 ] = fresh_wire_2026[ 7 ];
	assign fresh_wire_2045[ 8 ] = fresh_wire_2026[ 8 ];
	assign fresh_wire_2045[ 9 ] = fresh_wire_2026[ 9 ];
	assign fresh_wire_2045[ 10 ] = fresh_wire_2026[ 10 ];
	assign fresh_wire_2045[ 11 ] = fresh_wire_2026[ 11 ];
	assign fresh_wire_2045[ 12 ] = fresh_wire_2026[ 12 ];
	assign fresh_wire_2045[ 13 ] = fresh_wire_2026[ 13 ];
	assign fresh_wire_2045[ 14 ] = fresh_wire_2026[ 14 ];
	assign fresh_wire_2045[ 15 ] = fresh_wire_2026[ 15 ];
	assign fresh_wire_2047[ 0 ] = fresh_wire_2004[ 0 ];
	assign fresh_wire_2064[ 0 ] = fresh_wire_2068[ 0 ];
	assign fresh_wire_2064[ 1 ] = fresh_wire_2069[ 0 ];
	assign fresh_wire_2064[ 2 ] = fresh_wire_2070[ 0 ];
	assign fresh_wire_2064[ 3 ] = fresh_wire_2071[ 0 ];
	assign fresh_wire_2064[ 4 ] = fresh_wire_2072[ 0 ];
	assign fresh_wire_2064[ 5 ] = fresh_wire_2073[ 0 ];
	assign fresh_wire_2064[ 6 ] = fresh_wire_2074[ 0 ];
	assign fresh_wire_2064[ 7 ] = fresh_wire_2075[ 0 ];
	assign fresh_wire_2064[ 8 ] = fresh_wire_2076[ 0 ];
	assign fresh_wire_2065[ 0 ] = fresh_wire_1407[ 0 ];
	assign fresh_wire_2065[ 1 ] = fresh_wire_1407[ 1 ];
	assign fresh_wire_2065[ 2 ] = fresh_wire_1407[ 2 ];
	assign fresh_wire_2065[ 3 ] = fresh_wire_1407[ 3 ];
	assign fresh_wire_2065[ 4 ] = fresh_wire_1407[ 4 ];
	assign fresh_wire_2065[ 5 ] = fresh_wire_1407[ 5 ];
	assign fresh_wire_2065[ 6 ] = fresh_wire_1407[ 6 ];
	assign fresh_wire_2065[ 7 ] = fresh_wire_1407[ 7 ];
	assign fresh_wire_2065[ 8 ] = fresh_wire_1407[ 8 ];
	assign fresh_wire_2067[ 0 ] = fresh_wire_2007[ 0 ];
	assign fresh_wire_2077[ 0 ] = fresh_wire_2081[ 0 ];
	assign fresh_wire_2077[ 1 ] = fresh_wire_2082[ 0 ];
	assign fresh_wire_2077[ 2 ] = fresh_wire_2083[ 0 ];
	assign fresh_wire_2077[ 3 ] = fresh_wire_2084[ 0 ];
	assign fresh_wire_2077[ 4 ] = fresh_wire_2085[ 0 ];
	assign fresh_wire_2077[ 5 ] = fresh_wire_2086[ 0 ];
	assign fresh_wire_2077[ 6 ] = fresh_wire_2087[ 0 ];
	assign fresh_wire_2077[ 7 ] = fresh_wire_2088[ 0 ];
	assign fresh_wire_2077[ 8 ] = fresh_wire_2089[ 0 ];
	assign fresh_wire_2078[ 0 ] = fresh_wire_2066[ 0 ];
	assign fresh_wire_2078[ 1 ] = fresh_wire_2066[ 1 ];
	assign fresh_wire_2078[ 2 ] = fresh_wire_2066[ 2 ];
	assign fresh_wire_2078[ 3 ] = fresh_wire_2066[ 3 ];
	assign fresh_wire_2078[ 4 ] = fresh_wire_2066[ 4 ];
	assign fresh_wire_2078[ 5 ] = fresh_wire_2066[ 5 ];
	assign fresh_wire_2078[ 6 ] = fresh_wire_2066[ 6 ];
	assign fresh_wire_2078[ 7 ] = fresh_wire_2066[ 7 ];
	assign fresh_wire_2078[ 8 ] = fresh_wire_2066[ 8 ];
	assign fresh_wire_2080[ 0 ] = fresh_wire_2004[ 0 ];
	assign fresh_wire_2090[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_2091[ 0 ] = fresh_wire_1407[ 0 ];
	assign fresh_wire_2091[ 1 ] = fresh_wire_1407[ 1 ];
	assign fresh_wire_2091[ 2 ] = fresh_wire_1407[ 2 ];
	assign fresh_wire_2091[ 3 ] = fresh_wire_1407[ 3 ];
	assign fresh_wire_2091[ 4 ] = fresh_wire_1407[ 4 ];
	assign fresh_wire_2091[ 5 ] = fresh_wire_1407[ 5 ];
	assign fresh_wire_2091[ 6 ] = fresh_wire_1407[ 6 ];
	assign fresh_wire_2091[ 7 ] = fresh_wire_1407[ 7 ];
	assign fresh_wire_2091[ 8 ] = fresh_wire_1407[ 8 ];
	assign fresh_wire_2093[ 0 ] = fresh_wire_2079[ 0 ];
	assign fresh_wire_2093[ 1 ] = fresh_wire_2079[ 1 ];
	assign fresh_wire_2093[ 2 ] = fresh_wire_2079[ 2 ];
	assign fresh_wire_2093[ 3 ] = fresh_wire_2079[ 3 ];
	assign fresh_wire_2093[ 4 ] = fresh_wire_2079[ 4 ];
	assign fresh_wire_2093[ 5 ] = fresh_wire_2079[ 5 ];
	assign fresh_wire_2093[ 6 ] = fresh_wire_2079[ 6 ];
	assign fresh_wire_2093[ 7 ] = fresh_wire_2079[ 7 ];
	assign fresh_wire_2093[ 8 ] = fresh_wire_2079[ 8 ];
	assign fresh_wire_2094[ 0 ] = fresh_wire_2046[ 0 ];
	assign fresh_wire_2094[ 1 ] = fresh_wire_2046[ 1 ];
	assign fresh_wire_2094[ 2 ] = fresh_wire_2046[ 2 ];
	assign fresh_wire_2094[ 3 ] = fresh_wire_2046[ 3 ];
	assign fresh_wire_2094[ 4 ] = fresh_wire_2046[ 4 ];
	assign fresh_wire_2094[ 5 ] = fresh_wire_2046[ 5 ];
	assign fresh_wire_2094[ 6 ] = fresh_wire_2046[ 6 ];
	assign fresh_wire_2094[ 7 ] = fresh_wire_2046[ 7 ];
	assign fresh_wire_2094[ 8 ] = fresh_wire_2046[ 8 ];
	assign fresh_wire_2094[ 9 ] = fresh_wire_2046[ 9 ];
	assign fresh_wire_2094[ 10 ] = fresh_wire_2046[ 10 ];
	assign fresh_wire_2094[ 11 ] = fresh_wire_2046[ 11 ];
	assign fresh_wire_2094[ 12 ] = fresh_wire_2046[ 12 ];
	assign fresh_wire_2094[ 13 ] = fresh_wire_2046[ 13 ];
	assign fresh_wire_2094[ 14 ] = fresh_wire_2046[ 14 ];
	assign fresh_wire_2094[ 15 ] = fresh_wire_2046[ 15 ];
	assign fresh_wire_2095[ 0 ] = fresh_wire_2022[ 0 ];
	assign fresh_wire_2096[ 0 ] = fresh_wire_1581[ 0 ];
	assign fresh_wire_2096[ 1 ] = fresh_wire_1581[ 1 ];
	assign fresh_wire_2096[ 2 ] = fresh_wire_1581[ 2 ];
	assign fresh_wire_2096[ 3 ] = fresh_wire_1581[ 3 ];
	assign fresh_wire_2096[ 4 ] = fresh_wire_1581[ 4 ];
	assign fresh_wire_2096[ 5 ] = fresh_wire_1581[ 5 ];
	assign fresh_wire_2096[ 6 ] = fresh_wire_1581[ 6 ];
	assign fresh_wire_2096[ 7 ] = fresh_wire_1581[ 7 ];
	assign fresh_wire_2096[ 8 ] = fresh_wire_1581[ 8 ];
	assign fresh_wire_2096[ 9 ] = fresh_wire_1581[ 9 ];
	assign fresh_wire_2096[ 10 ] = fresh_wire_1581[ 10 ];
	assign fresh_wire_2096[ 11 ] = fresh_wire_1581[ 11 ];
	assign fresh_wire_2096[ 12 ] = fresh_wire_1581[ 12 ];
	assign fresh_wire_2096[ 13 ] = fresh_wire_1581[ 13 ];
	assign fresh_wire_2096[ 14 ] = fresh_wire_1581[ 14 ];
	assign fresh_wire_2096[ 15 ] = fresh_wire_1581[ 15 ];
	assign fresh_wire_2098[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_2099[ 0 ] = fresh_wire_96[ 0 ];
	assign fresh_wire_2099[ 1 ] = fresh_wire_94[ 0 ];
	assign fresh_wire_2099[ 2 ] = fresh_wire_92[ 0 ];
	assign fresh_wire_2099[ 3 ] = fresh_wire_90[ 0 ];
	assign fresh_wire_2099[ 4 ] = fresh_wire_88[ 0 ];
	assign fresh_wire_2099[ 5 ] = fresh_wire_86[ 0 ];
	assign fresh_wire_2099[ 6 ] = fresh_wire_114[ 0 ];
	assign fresh_wire_2099[ 7 ] = fresh_wire_112[ 0 ];
	assign fresh_wire_2099[ 8 ] = fresh_wire_110[ 0 ];
	assign fresh_wire_2099[ 9 ] = fresh_wire_108[ 0 ];
	assign fresh_wire_2099[ 10 ] = fresh_wire_106[ 0 ];
	assign fresh_wire_2099[ 11 ] = fresh_wire_104[ 0 ];
	assign fresh_wire_2099[ 12 ] = fresh_wire_102[ 0 ];
	assign fresh_wire_2099[ 13 ] = fresh_wire_100[ 0 ];
	assign fresh_wire_2099[ 14 ] = fresh_wire_98[ 0 ];
	assign fresh_wire_2099[ 15 ] = fresh_wire_84[ 0 ];
	assign fresh_wire_2101[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_2102[ 0 ] = fresh_wire_96[ 0 ];
	assign fresh_wire_2102[ 1 ] = fresh_wire_94[ 0 ];
	assign fresh_wire_2102[ 2 ] = fresh_wire_92[ 0 ];
	assign fresh_wire_2102[ 3 ] = fresh_wire_90[ 0 ];
	assign fresh_wire_2102[ 4 ] = fresh_wire_88[ 0 ];
	assign fresh_wire_2102[ 5 ] = fresh_wire_86[ 0 ];
	assign fresh_wire_2102[ 6 ] = fresh_wire_114[ 0 ];
	assign fresh_wire_2102[ 7 ] = fresh_wire_112[ 0 ];
	assign fresh_wire_2102[ 8 ] = fresh_wire_110[ 0 ];
	assign fresh_wire_2102[ 9 ] = fresh_wire_108[ 0 ];
	assign fresh_wire_2102[ 10 ] = fresh_wire_106[ 0 ];
	assign fresh_wire_2102[ 11 ] = fresh_wire_104[ 0 ];
	assign fresh_wire_2102[ 12 ] = fresh_wire_102[ 0 ];
	assign fresh_wire_2102[ 13 ] = fresh_wire_100[ 0 ];
	assign fresh_wire_2102[ 14 ] = fresh_wire_98[ 0 ];
	assign fresh_wire_2102[ 15 ] = fresh_wire_84[ 0 ];
	assign fresh_wire_2102[ 16 ] = fresh_wire_2269[ 0 ];
	assign fresh_wire_2104[ 0 ] = fresh_wire_2103[ 0 ];
	assign fresh_wire_2104[ 1 ] = fresh_wire_2103[ 1 ];
	assign fresh_wire_2104[ 2 ] = fresh_wire_2103[ 2 ];
	assign fresh_wire_2104[ 3 ] = fresh_wire_2103[ 3 ];
	assign fresh_wire_2104[ 4 ] = fresh_wire_2103[ 4 ];
	assign fresh_wire_2104[ 5 ] = fresh_wire_2103[ 5 ];
	assign fresh_wire_2104[ 6 ] = fresh_wire_2103[ 6 ];
	assign fresh_wire_2104[ 7 ] = fresh_wire_2103[ 7 ];
	assign fresh_wire_2104[ 8 ] = fresh_wire_2103[ 8 ];
	assign fresh_wire_2104[ 9 ] = fresh_wire_2103[ 9 ];
	assign fresh_wire_2104[ 10 ] = fresh_wire_2103[ 10 ];
	assign fresh_wire_2104[ 11 ] = fresh_wire_2103[ 11 ];
	assign fresh_wire_2104[ 12 ] = fresh_wire_2103[ 12 ];
	assign fresh_wire_2104[ 13 ] = fresh_wire_2103[ 13 ];
	assign fresh_wire_2104[ 14 ] = fresh_wire_2103[ 14 ];
	assign fresh_wire_2104[ 15 ] = fresh_wire_2103[ 15 ];
	assign fresh_wire_2104[ 16 ] = fresh_wire_2103[ 16 ];
	assign fresh_wire_2104[ 17 ] = fresh_wire_2103[ 17 ];
	assign fresh_wire_2104[ 18 ] = fresh_wire_2103[ 18 ];
	assign fresh_wire_2104[ 19 ] = fresh_wire_2103[ 19 ];
	assign fresh_wire_2104[ 20 ] = fresh_wire_2103[ 20 ];
	assign fresh_wire_2104[ 21 ] = fresh_wire_2103[ 21 ];
	assign fresh_wire_2104[ 22 ] = fresh_wire_2103[ 22 ];
	assign fresh_wire_2104[ 23 ] = fresh_wire_2103[ 23 ];
	assign fresh_wire_2104[ 24 ] = fresh_wire_2103[ 24 ];
	assign fresh_wire_2104[ 25 ] = fresh_wire_2103[ 25 ];
	assign fresh_wire_2104[ 26 ] = fresh_wire_2103[ 26 ];
	assign fresh_wire_2104[ 27 ] = fresh_wire_2103[ 27 ];
	assign fresh_wire_2104[ 28 ] = fresh_wire_2103[ 28 ];
	assign fresh_wire_2104[ 29 ] = fresh_wire_2103[ 29 ];
	assign fresh_wire_2104[ 30 ] = fresh_wire_2103[ 30 ];
	assign fresh_wire_2104[ 31 ] = fresh_wire_2103[ 31 ];
	assign fresh_wire_2104[ 32 ] = fresh_wire_2103[ 32 ];
	assign fresh_wire_2104[ 33 ] = fresh_wire_2103[ 33 ];
	assign fresh_wire_2105[ 0 ] = fresh_wire_2270[ 0 ];
	assign fresh_wire_2105[ 1 ] = fresh_wire_2270[ 1 ];
	assign fresh_wire_2105[ 2 ] = fresh_wire_2270[ 2 ];
	assign fresh_wire_2105[ 3 ] = fresh_wire_2270[ 3 ];
	assign fresh_wire_2105[ 4 ] = fresh_wire_2270[ 4 ];
	assign fresh_wire_2105[ 5 ] = fresh_wire_2270[ 5 ];
	assign fresh_wire_2105[ 6 ] = fresh_wire_2270[ 6 ];
	assign fresh_wire_2105[ 7 ] = fresh_wire_2270[ 7 ];
	assign fresh_wire_2105[ 8 ] = fresh_wire_2270[ 8 ];
	assign fresh_wire_2105[ 9 ] = fresh_wire_2270[ 9 ];
	assign fresh_wire_2105[ 10 ] = fresh_wire_2270[ 10 ];
	assign fresh_wire_2105[ 11 ] = fresh_wire_2270[ 11 ];
	assign fresh_wire_2105[ 12 ] = fresh_wire_2270[ 12 ];
	assign fresh_wire_2105[ 13 ] = fresh_wire_2270[ 13 ];
	assign fresh_wire_2105[ 14 ] = fresh_wire_2270[ 14 ];
	assign fresh_wire_2105[ 15 ] = fresh_wire_2270[ 15 ];
	assign fresh_wire_2105[ 16 ] = fresh_wire_2270[ 16 ];
	assign fresh_wire_2105[ 17 ] = fresh_wire_2270[ 17 ];
	assign fresh_wire_2105[ 18 ] = fresh_wire_2270[ 18 ];
	assign fresh_wire_2105[ 19 ] = fresh_wire_2270[ 19 ];
	assign fresh_wire_2105[ 20 ] = fresh_wire_2270[ 20 ];
	assign fresh_wire_2105[ 21 ] = fresh_wire_2270[ 21 ];
	assign fresh_wire_2105[ 22 ] = fresh_wire_2270[ 22 ];
	assign fresh_wire_2105[ 23 ] = fresh_wire_2270[ 23 ];
	assign fresh_wire_2105[ 24 ] = fresh_wire_2270[ 24 ];
	assign fresh_wire_2105[ 25 ] = fresh_wire_2270[ 25 ];
	assign fresh_wire_2105[ 26 ] = fresh_wire_2270[ 26 ];
	assign fresh_wire_2105[ 27 ] = fresh_wire_2270[ 27 ];
	assign fresh_wire_2105[ 28 ] = fresh_wire_2270[ 28 ];
	assign fresh_wire_2105[ 29 ] = fresh_wire_2270[ 29 ];
	assign fresh_wire_2105[ 30 ] = fresh_wire_2270[ 30 ];
	assign fresh_wire_2105[ 31 ] = fresh_wire_2270[ 31 ];
	assign fresh_wire_2105[ 32 ] = fresh_wire_2270[ 32 ];
	assign fresh_wire_2105[ 33 ] = fresh_wire_2270[ 33 ];
	assign fresh_wire_2107[ 0 ] = fresh_wire_2100[ 0 ];
	assign fresh_wire_2107[ 1 ] = fresh_wire_2100[ 1 ];
	assign fresh_wire_2107[ 2 ] = fresh_wire_2100[ 2 ];
	assign fresh_wire_2107[ 3 ] = fresh_wire_2100[ 3 ];
	assign fresh_wire_2107[ 4 ] = fresh_wire_2100[ 4 ];
	assign fresh_wire_2107[ 5 ] = fresh_wire_2100[ 5 ];
	assign fresh_wire_2107[ 6 ] = fresh_wire_2100[ 6 ];
	assign fresh_wire_2107[ 7 ] = fresh_wire_2100[ 7 ];
	assign fresh_wire_2107[ 8 ] = fresh_wire_2100[ 8 ];
	assign fresh_wire_2107[ 9 ] = fresh_wire_2100[ 9 ];
	assign fresh_wire_2107[ 10 ] = fresh_wire_2100[ 10 ];
	assign fresh_wire_2107[ 11 ] = fresh_wire_2100[ 11 ];
	assign fresh_wire_2107[ 12 ] = fresh_wire_2100[ 12 ];
	assign fresh_wire_2107[ 13 ] = fresh_wire_2100[ 13 ];
	assign fresh_wire_2107[ 14 ] = fresh_wire_2100[ 14 ];
	assign fresh_wire_2107[ 15 ] = fresh_wire_2100[ 15 ];
	assign fresh_wire_2107[ 16 ] = fresh_wire_2271[ 0 ];
	assign fresh_wire_2109[ 0 ] = fresh_wire_2108[ 0 ];
	assign fresh_wire_2109[ 1 ] = fresh_wire_2108[ 1 ];
	assign fresh_wire_2109[ 2 ] = fresh_wire_2108[ 2 ];
	assign fresh_wire_2109[ 3 ] = fresh_wire_2108[ 3 ];
	assign fresh_wire_2109[ 4 ] = fresh_wire_2108[ 4 ];
	assign fresh_wire_2109[ 5 ] = fresh_wire_2108[ 5 ];
	assign fresh_wire_2109[ 6 ] = fresh_wire_2108[ 6 ];
	assign fresh_wire_2109[ 7 ] = fresh_wire_2108[ 7 ];
	assign fresh_wire_2109[ 8 ] = fresh_wire_2108[ 8 ];
	assign fresh_wire_2109[ 9 ] = fresh_wire_2108[ 9 ];
	assign fresh_wire_2109[ 10 ] = fresh_wire_2108[ 10 ];
	assign fresh_wire_2109[ 11 ] = fresh_wire_2108[ 11 ];
	assign fresh_wire_2109[ 12 ] = fresh_wire_2108[ 12 ];
	assign fresh_wire_2109[ 13 ] = fresh_wire_2108[ 13 ];
	assign fresh_wire_2109[ 14 ] = fresh_wire_2108[ 14 ];
	assign fresh_wire_2109[ 15 ] = fresh_wire_2108[ 15 ];
	assign fresh_wire_2109[ 16 ] = fresh_wire_2108[ 16 ];
	assign fresh_wire_2109[ 17 ] = fresh_wire_2108[ 17 ];
	assign fresh_wire_2109[ 18 ] = fresh_wire_2108[ 18 ];
	assign fresh_wire_2109[ 19 ] = fresh_wire_2108[ 19 ];
	assign fresh_wire_2109[ 20 ] = fresh_wire_2108[ 20 ];
	assign fresh_wire_2109[ 21 ] = fresh_wire_2108[ 21 ];
	assign fresh_wire_2109[ 22 ] = fresh_wire_2108[ 22 ];
	assign fresh_wire_2109[ 23 ] = fresh_wire_2108[ 23 ];
	assign fresh_wire_2109[ 24 ] = fresh_wire_2108[ 24 ];
	assign fresh_wire_2109[ 25 ] = fresh_wire_2108[ 25 ];
	assign fresh_wire_2109[ 26 ] = fresh_wire_2108[ 26 ];
	assign fresh_wire_2109[ 27 ] = fresh_wire_2108[ 27 ];
	assign fresh_wire_2109[ 28 ] = fresh_wire_2108[ 28 ];
	assign fresh_wire_2109[ 29 ] = fresh_wire_2108[ 29 ];
	assign fresh_wire_2109[ 30 ] = fresh_wire_2108[ 30 ];
	assign fresh_wire_2109[ 31 ] = fresh_wire_2108[ 31 ];
	assign fresh_wire_2109[ 32 ] = fresh_wire_2108[ 32 ];
	assign fresh_wire_2109[ 33 ] = fresh_wire_2108[ 33 ];
	assign fresh_wire_2110[ 0 ] = fresh_wire_2272[ 0 ];
	assign fresh_wire_2110[ 1 ] = fresh_wire_2272[ 1 ];
	assign fresh_wire_2110[ 2 ] = fresh_wire_2272[ 2 ];
	assign fresh_wire_2110[ 3 ] = fresh_wire_2272[ 3 ];
	assign fresh_wire_2110[ 4 ] = fresh_wire_2272[ 4 ];
	assign fresh_wire_2110[ 5 ] = fresh_wire_2272[ 5 ];
	assign fresh_wire_2110[ 6 ] = fresh_wire_2272[ 6 ];
	assign fresh_wire_2110[ 7 ] = fresh_wire_2272[ 7 ];
	assign fresh_wire_2110[ 8 ] = fresh_wire_2272[ 8 ];
	assign fresh_wire_2110[ 9 ] = fresh_wire_2272[ 9 ];
	assign fresh_wire_2110[ 10 ] = fresh_wire_2272[ 10 ];
	assign fresh_wire_2110[ 11 ] = fresh_wire_2272[ 11 ];
	assign fresh_wire_2110[ 12 ] = fresh_wire_2272[ 12 ];
	assign fresh_wire_2110[ 13 ] = fresh_wire_2272[ 13 ];
	assign fresh_wire_2110[ 14 ] = fresh_wire_2272[ 14 ];
	assign fresh_wire_2110[ 15 ] = fresh_wire_2272[ 15 ];
	assign fresh_wire_2110[ 16 ] = fresh_wire_2272[ 16 ];
	assign fresh_wire_2110[ 17 ] = fresh_wire_2272[ 17 ];
	assign fresh_wire_2110[ 18 ] = fresh_wire_2272[ 18 ];
	assign fresh_wire_2110[ 19 ] = fresh_wire_2272[ 19 ];
	assign fresh_wire_2110[ 20 ] = fresh_wire_2272[ 20 ];
	assign fresh_wire_2110[ 21 ] = fresh_wire_2272[ 21 ];
	assign fresh_wire_2110[ 22 ] = fresh_wire_2272[ 22 ];
	assign fresh_wire_2110[ 23 ] = fresh_wire_2272[ 23 ];
	assign fresh_wire_2110[ 24 ] = fresh_wire_2272[ 24 ];
	assign fresh_wire_2110[ 25 ] = fresh_wire_2272[ 25 ];
	assign fresh_wire_2110[ 26 ] = fresh_wire_2272[ 26 ];
	assign fresh_wire_2110[ 27 ] = fresh_wire_2272[ 27 ];
	assign fresh_wire_2110[ 28 ] = fresh_wire_2272[ 28 ];
	assign fresh_wire_2110[ 29 ] = fresh_wire_2272[ 29 ];
	assign fresh_wire_2110[ 30 ] = fresh_wire_2272[ 30 ];
	assign fresh_wire_2110[ 31 ] = fresh_wire_2272[ 31 ];
	assign fresh_wire_2110[ 32 ] = fresh_wire_2272[ 32 ];
	assign fresh_wire_2110[ 33 ] = fresh_wire_2272[ 33 ];
	assign fresh_wire_2112[ 0 ] = fresh_wire_609[ 0 ];
	assign fresh_wire_2112[ 1 ] = fresh_wire_609[ 1 ];
	assign fresh_wire_2112[ 2 ] = fresh_wire_609[ 2 ];
	assign fresh_wire_2112[ 3 ] = fresh_wire_609[ 3 ];
	assign fresh_wire_2112[ 4 ] = fresh_wire_609[ 4 ];
	assign fresh_wire_2112[ 5 ] = fresh_wire_609[ 5 ];
	assign fresh_wire_2112[ 6 ] = fresh_wire_609[ 6 ];
	assign fresh_wire_2112[ 7 ] = fresh_wire_609[ 7 ];
	assign fresh_wire_2112[ 8 ] = fresh_wire_609[ 8 ];
	assign fresh_wire_2112[ 9 ] = fresh_wire_609[ 9 ];
	assign fresh_wire_2112[ 10 ] = fresh_wire_609[ 10 ];
	assign fresh_wire_2112[ 11 ] = fresh_wire_609[ 11 ];
	assign fresh_wire_2112[ 12 ] = fresh_wire_609[ 12 ];
	assign fresh_wire_2112[ 13 ] = fresh_wire_609[ 13 ];
	assign fresh_wire_2112[ 14 ] = fresh_wire_609[ 14 ];
	assign fresh_wire_2112[ 15 ] = fresh_wire_609[ 15 ];
	assign fresh_wire_2112[ 16 ] = fresh_wire_2273[ 0 ];
	assign fresh_wire_2114[ 0 ] = fresh_wire_2113[ 0 ];
	assign fresh_wire_2114[ 1 ] = fresh_wire_2113[ 1 ];
	assign fresh_wire_2114[ 2 ] = fresh_wire_2113[ 2 ];
	assign fresh_wire_2114[ 3 ] = fresh_wire_2113[ 3 ];
	assign fresh_wire_2114[ 4 ] = fresh_wire_2113[ 4 ];
	assign fresh_wire_2114[ 5 ] = fresh_wire_2113[ 5 ];
	assign fresh_wire_2114[ 6 ] = fresh_wire_2113[ 6 ];
	assign fresh_wire_2114[ 7 ] = fresh_wire_2113[ 7 ];
	assign fresh_wire_2114[ 8 ] = fresh_wire_2113[ 8 ];
	assign fresh_wire_2114[ 9 ] = fresh_wire_2113[ 9 ];
	assign fresh_wire_2114[ 10 ] = fresh_wire_2113[ 10 ];
	assign fresh_wire_2114[ 11 ] = fresh_wire_2113[ 11 ];
	assign fresh_wire_2114[ 12 ] = fresh_wire_2113[ 12 ];
	assign fresh_wire_2114[ 13 ] = fresh_wire_2113[ 13 ];
	assign fresh_wire_2114[ 14 ] = fresh_wire_2113[ 14 ];
	assign fresh_wire_2114[ 15 ] = fresh_wire_2113[ 15 ];
	assign fresh_wire_2114[ 16 ] = fresh_wire_2113[ 16 ];
	assign fresh_wire_2114[ 17 ] = fresh_wire_2113[ 17 ];
	assign fresh_wire_2114[ 18 ] = fresh_wire_2113[ 18 ];
	assign fresh_wire_2114[ 19 ] = fresh_wire_2113[ 19 ];
	assign fresh_wire_2114[ 20 ] = fresh_wire_2113[ 20 ];
	assign fresh_wire_2114[ 21 ] = fresh_wire_2113[ 21 ];
	assign fresh_wire_2114[ 22 ] = fresh_wire_2113[ 22 ];
	assign fresh_wire_2114[ 23 ] = fresh_wire_2113[ 23 ];
	assign fresh_wire_2114[ 24 ] = fresh_wire_2113[ 24 ];
	assign fresh_wire_2114[ 25 ] = fresh_wire_2113[ 25 ];
	assign fresh_wire_2114[ 26 ] = fresh_wire_2113[ 26 ];
	assign fresh_wire_2114[ 27 ] = fresh_wire_2113[ 27 ];
	assign fresh_wire_2114[ 28 ] = fresh_wire_2113[ 28 ];
	assign fresh_wire_2114[ 29 ] = fresh_wire_2113[ 29 ];
	assign fresh_wire_2114[ 30 ] = fresh_wire_2113[ 30 ];
	assign fresh_wire_2114[ 31 ] = fresh_wire_2113[ 31 ];
	assign fresh_wire_2114[ 32 ] = fresh_wire_2113[ 32 ];
	assign fresh_wire_2114[ 33 ] = fresh_wire_2113[ 33 ];
	assign fresh_wire_2115[ 0 ] = fresh_wire_2274[ 0 ];
	assign fresh_wire_2115[ 1 ] = fresh_wire_2274[ 1 ];
	assign fresh_wire_2115[ 2 ] = fresh_wire_2274[ 2 ];
	assign fresh_wire_2115[ 3 ] = fresh_wire_2274[ 3 ];
	assign fresh_wire_2115[ 4 ] = fresh_wire_2274[ 4 ];
	assign fresh_wire_2115[ 5 ] = fresh_wire_2274[ 5 ];
	assign fresh_wire_2115[ 6 ] = fresh_wire_2274[ 6 ];
	assign fresh_wire_2115[ 7 ] = fresh_wire_2274[ 7 ];
	assign fresh_wire_2115[ 8 ] = fresh_wire_2274[ 8 ];
	assign fresh_wire_2115[ 9 ] = fresh_wire_2274[ 9 ];
	assign fresh_wire_2115[ 10 ] = fresh_wire_2274[ 10 ];
	assign fresh_wire_2115[ 11 ] = fresh_wire_2274[ 11 ];
	assign fresh_wire_2115[ 12 ] = fresh_wire_2274[ 12 ];
	assign fresh_wire_2115[ 13 ] = fresh_wire_2274[ 13 ];
	assign fresh_wire_2115[ 14 ] = fresh_wire_2274[ 14 ];
	assign fresh_wire_2115[ 15 ] = fresh_wire_2274[ 15 ];
	assign fresh_wire_2115[ 16 ] = fresh_wire_2274[ 16 ];
	assign fresh_wire_2115[ 17 ] = fresh_wire_2274[ 17 ];
	assign fresh_wire_2115[ 18 ] = fresh_wire_2274[ 18 ];
	assign fresh_wire_2115[ 19 ] = fresh_wire_2274[ 19 ];
	assign fresh_wire_2115[ 20 ] = fresh_wire_2274[ 20 ];
	assign fresh_wire_2115[ 21 ] = fresh_wire_2274[ 21 ];
	assign fresh_wire_2115[ 22 ] = fresh_wire_2274[ 22 ];
	assign fresh_wire_2115[ 23 ] = fresh_wire_2274[ 23 ];
	assign fresh_wire_2115[ 24 ] = fresh_wire_2274[ 24 ];
	assign fresh_wire_2115[ 25 ] = fresh_wire_2274[ 25 ];
	assign fresh_wire_2115[ 26 ] = fresh_wire_2274[ 26 ];
	assign fresh_wire_2115[ 27 ] = fresh_wire_2274[ 27 ];
	assign fresh_wire_2115[ 28 ] = fresh_wire_2274[ 28 ];
	assign fresh_wire_2115[ 29 ] = fresh_wire_2274[ 29 ];
	assign fresh_wire_2115[ 30 ] = fresh_wire_2274[ 30 ];
	assign fresh_wire_2115[ 31 ] = fresh_wire_2274[ 31 ];
	assign fresh_wire_2115[ 32 ] = fresh_wire_2274[ 32 ];
	assign fresh_wire_2115[ 33 ] = fresh_wire_2274[ 33 ];
	assign fresh_wire_2118[ 0 ] = fresh_wire_2137[ 0 ];
	assign fresh_wire_2118[ 1 ] = fresh_wire_2137[ 1 ];
	assign fresh_wire_2118[ 2 ] = fresh_wire_2137[ 2 ];
	assign fresh_wire_2118[ 3 ] = fresh_wire_2137[ 3 ];
	assign fresh_wire_2118[ 4 ] = fresh_wire_2137[ 4 ];
	assign fresh_wire_2118[ 5 ] = fresh_wire_2137[ 5 ];
	assign fresh_wire_2118[ 6 ] = fresh_wire_2137[ 6 ];
	assign fresh_wire_2118[ 7 ] = fresh_wire_2137[ 7 ];
	assign fresh_wire_2118[ 8 ] = fresh_wire_2137[ 8 ];
	assign fresh_wire_2118[ 9 ] = fresh_wire_2137[ 9 ];
	assign fresh_wire_2118[ 10 ] = fresh_wire_2137[ 10 ];
	assign fresh_wire_2118[ 11 ] = fresh_wire_2137[ 11 ];
	assign fresh_wire_2118[ 12 ] = fresh_wire_2137[ 12 ];
	assign fresh_wire_2118[ 13 ] = fresh_wire_2137[ 13 ];
	assign fresh_wire_2118[ 14 ] = fresh_wire_2137[ 14 ];
	assign fresh_wire_2118[ 15 ] = fresh_wire_2137[ 15 ];
	assign fresh_wire_2120[ 0 ] = fresh_wire_2142[ 0 ];
	assign fresh_wire_2120[ 1 ] = fresh_wire_2142[ 1 ];
	assign fresh_wire_2120[ 2 ] = fresh_wire_2142[ 2 ];
	assign fresh_wire_2120[ 3 ] = fresh_wire_2142[ 3 ];
	assign fresh_wire_2120[ 4 ] = fresh_wire_2142[ 4 ];
	assign fresh_wire_2120[ 5 ] = fresh_wire_2142[ 5 ];
	assign fresh_wire_2120[ 6 ] = fresh_wire_2142[ 6 ];
	assign fresh_wire_2120[ 7 ] = fresh_wire_2142[ 7 ];
	assign fresh_wire_2120[ 8 ] = fresh_wire_2142[ 8 ];
	assign fresh_wire_2120[ 9 ] = fresh_wire_2142[ 9 ];
	assign fresh_wire_2120[ 10 ] = fresh_wire_2142[ 10 ];
	assign fresh_wire_2120[ 11 ] = fresh_wire_2142[ 11 ];
	assign fresh_wire_2120[ 12 ] = fresh_wire_2142[ 12 ];
	assign fresh_wire_2120[ 13 ] = fresh_wire_2142[ 13 ];
	assign fresh_wire_2120[ 14 ] = fresh_wire_2142[ 14 ];
	assign fresh_wire_2120[ 15 ] = fresh_wire_2142[ 15 ];
	assign fresh_wire_2122[ 0 ] = fresh_wire_2119[ 0 ];
	assign fresh_wire_2122[ 1 ] = fresh_wire_2119[ 1 ];
	assign fresh_wire_2122[ 2 ] = fresh_wire_2119[ 2 ];
	assign fresh_wire_2122[ 3 ] = fresh_wire_2119[ 3 ];
	assign fresh_wire_2122[ 4 ] = fresh_wire_2119[ 4 ];
	assign fresh_wire_2122[ 5 ] = fresh_wire_2119[ 5 ];
	assign fresh_wire_2122[ 6 ] = fresh_wire_2119[ 6 ];
	assign fresh_wire_2122[ 7 ] = fresh_wire_2119[ 7 ];
	assign fresh_wire_2122[ 8 ] = fresh_wire_2119[ 8 ];
	assign fresh_wire_2122[ 9 ] = fresh_wire_2119[ 9 ];
	assign fresh_wire_2122[ 10 ] = fresh_wire_2119[ 10 ];
	assign fresh_wire_2122[ 11 ] = fresh_wire_2119[ 11 ];
	assign fresh_wire_2122[ 12 ] = fresh_wire_2119[ 12 ];
	assign fresh_wire_2122[ 13 ] = fresh_wire_2119[ 13 ];
	assign fresh_wire_2122[ 14 ] = fresh_wire_2119[ 14 ];
	assign fresh_wire_2122[ 15 ] = fresh_wire_2119[ 15 ];
	assign fresh_wire_2122[ 16 ] = fresh_wire_2119[ 16 ];
	assign fresh_wire_2123[ 0 ] = fresh_wire_2121[ 0 ];
	assign fresh_wire_2123[ 1 ] = fresh_wire_2121[ 1 ];
	assign fresh_wire_2123[ 2 ] = fresh_wire_2121[ 2 ];
	assign fresh_wire_2123[ 3 ] = fresh_wire_2121[ 3 ];
	assign fresh_wire_2123[ 4 ] = fresh_wire_2121[ 4 ];
	assign fresh_wire_2123[ 5 ] = fresh_wire_2121[ 5 ];
	assign fresh_wire_2123[ 6 ] = fresh_wire_2121[ 6 ];
	assign fresh_wire_2123[ 7 ] = fresh_wire_2121[ 7 ];
	assign fresh_wire_2123[ 8 ] = fresh_wire_2121[ 8 ];
	assign fresh_wire_2123[ 9 ] = fresh_wire_2121[ 9 ];
	assign fresh_wire_2123[ 10 ] = fresh_wire_2121[ 10 ];
	assign fresh_wire_2123[ 11 ] = fresh_wire_2121[ 11 ];
	assign fresh_wire_2123[ 12 ] = fresh_wire_2121[ 12 ];
	assign fresh_wire_2123[ 13 ] = fresh_wire_2121[ 13 ];
	assign fresh_wire_2123[ 14 ] = fresh_wire_2121[ 14 ];
	assign fresh_wire_2123[ 15 ] = fresh_wire_2121[ 15 ];
	assign fresh_wire_2123[ 16 ] = fresh_wire_2121[ 16 ];
	assign fresh_wire_2125[ 0 ] = fresh_wire_2124[ 0 ];
	assign fresh_wire_2125[ 1 ] = fresh_wire_2124[ 1 ];
	assign fresh_wire_2125[ 2 ] = fresh_wire_2124[ 2 ];
	assign fresh_wire_2125[ 3 ] = fresh_wire_2124[ 3 ];
	assign fresh_wire_2125[ 4 ] = fresh_wire_2124[ 4 ];
	assign fresh_wire_2125[ 5 ] = fresh_wire_2124[ 5 ];
	assign fresh_wire_2125[ 6 ] = fresh_wire_2124[ 6 ];
	assign fresh_wire_2125[ 7 ] = fresh_wire_2124[ 7 ];
	assign fresh_wire_2125[ 8 ] = fresh_wire_2124[ 8 ];
	assign fresh_wire_2125[ 9 ] = fresh_wire_2124[ 9 ];
	assign fresh_wire_2125[ 10 ] = fresh_wire_2124[ 10 ];
	assign fresh_wire_2125[ 11 ] = fresh_wire_2124[ 11 ];
	assign fresh_wire_2125[ 12 ] = fresh_wire_2124[ 12 ];
	assign fresh_wire_2125[ 13 ] = fresh_wire_2124[ 13 ];
	assign fresh_wire_2125[ 14 ] = fresh_wire_2124[ 14 ];
	assign fresh_wire_2125[ 15 ] = fresh_wire_2124[ 15 ];
	assign fresh_wire_2125[ 16 ] = fresh_wire_2124[ 16 ];
	assign fresh_wire_2126[ 0 ] = fresh_wire_2279[ 0 ];
	assign fresh_wire_2126[ 1 ] = fresh_wire_2279[ 1 ];
	assign fresh_wire_2126[ 2 ] = fresh_wire_2279[ 2 ];
	assign fresh_wire_2126[ 3 ] = fresh_wire_2279[ 3 ];
	assign fresh_wire_2126[ 4 ] = fresh_wire_2279[ 4 ];
	assign fresh_wire_2126[ 5 ] = fresh_wire_2279[ 5 ];
	assign fresh_wire_2126[ 6 ] = fresh_wire_2279[ 6 ];
	assign fresh_wire_2126[ 7 ] = fresh_wire_2279[ 7 ];
	assign fresh_wire_2126[ 8 ] = fresh_wire_2279[ 8 ];
	assign fresh_wire_2126[ 9 ] = fresh_wire_2279[ 9 ];
	assign fresh_wire_2126[ 10 ] = fresh_wire_2279[ 10 ];
	assign fresh_wire_2126[ 11 ] = fresh_wire_2279[ 11 ];
	assign fresh_wire_2126[ 12 ] = fresh_wire_2279[ 12 ];
	assign fresh_wire_2126[ 13 ] = fresh_wire_2279[ 13 ];
	assign fresh_wire_2126[ 14 ] = fresh_wire_2279[ 14 ];
	assign fresh_wire_2126[ 15 ] = fresh_wire_2279[ 15 ];
	assign fresh_wire_2126[ 16 ] = fresh_wire_2279[ 16 ];
	assign fresh_wire_2128[ 0 ] = fresh_wire_2171[ 0 ];
	assign fresh_wire_2128[ 1 ] = fresh_wire_2171[ 1 ];
	assign fresh_wire_2128[ 2 ] = fresh_wire_2171[ 2 ];
	assign fresh_wire_2128[ 3 ] = fresh_wire_2171[ 3 ];
	assign fresh_wire_2128[ 4 ] = fresh_wire_2171[ 4 ];
	assign fresh_wire_2128[ 5 ] = fresh_wire_2171[ 5 ];
	assign fresh_wire_2128[ 6 ] = fresh_wire_2171[ 6 ];
	assign fresh_wire_2128[ 7 ] = fresh_wire_2171[ 7 ];
	assign fresh_wire_2128[ 8 ] = fresh_wire_2171[ 8 ];
	assign fresh_wire_2128[ 9 ] = fresh_wire_2171[ 9 ];
	assign fresh_wire_2128[ 10 ] = fresh_wire_2171[ 10 ];
	assign fresh_wire_2128[ 11 ] = fresh_wire_2171[ 11 ];
	assign fresh_wire_2128[ 12 ] = fresh_wire_2171[ 12 ];
	assign fresh_wire_2128[ 13 ] = fresh_wire_2171[ 13 ];
	assign fresh_wire_2128[ 14 ] = fresh_wire_2171[ 14 ];
	assign fresh_wire_2128[ 15 ] = fresh_wire_2171[ 15 ];
	assign fresh_wire_2130[ 0 ] = fresh_wire_2151[ 0 ];
	assign fresh_wire_2130[ 1 ] = fresh_wire_2151[ 1 ];
	assign fresh_wire_2130[ 2 ] = fresh_wire_2151[ 2 ];
	assign fresh_wire_2130[ 3 ] = fresh_wire_2151[ 3 ];
	assign fresh_wire_2130[ 4 ] = fresh_wire_2151[ 4 ];
	assign fresh_wire_2130[ 5 ] = fresh_wire_2151[ 5 ];
	assign fresh_wire_2130[ 6 ] = fresh_wire_2151[ 6 ];
	assign fresh_wire_2130[ 7 ] = fresh_wire_2151[ 7 ];
	assign fresh_wire_2130[ 8 ] = fresh_wire_2151[ 8 ];
	assign fresh_wire_2130[ 9 ] = fresh_wire_2151[ 9 ];
	assign fresh_wire_2130[ 10 ] = fresh_wire_2151[ 10 ];
	assign fresh_wire_2130[ 11 ] = fresh_wire_2151[ 11 ];
	assign fresh_wire_2130[ 12 ] = fresh_wire_2151[ 12 ];
	assign fresh_wire_2130[ 13 ] = fresh_wire_2151[ 13 ];
	assign fresh_wire_2130[ 14 ] = fresh_wire_2151[ 14 ];
	assign fresh_wire_2130[ 15 ] = fresh_wire_2151[ 15 ];
	assign fresh_wire_2132[ 0 ] = fresh_wire_2129[ 0 ];
	assign fresh_wire_2132[ 1 ] = fresh_wire_2129[ 1 ];
	assign fresh_wire_2132[ 2 ] = fresh_wire_2129[ 2 ];
	assign fresh_wire_2132[ 3 ] = fresh_wire_2129[ 3 ];
	assign fresh_wire_2132[ 4 ] = fresh_wire_2129[ 4 ];
	assign fresh_wire_2132[ 5 ] = fresh_wire_2129[ 5 ];
	assign fresh_wire_2132[ 6 ] = fresh_wire_2129[ 6 ];
	assign fresh_wire_2132[ 7 ] = fresh_wire_2129[ 7 ];
	assign fresh_wire_2132[ 8 ] = fresh_wire_2129[ 8 ];
	assign fresh_wire_2132[ 9 ] = fresh_wire_2129[ 9 ];
	assign fresh_wire_2132[ 10 ] = fresh_wire_2129[ 10 ];
	assign fresh_wire_2132[ 11 ] = fresh_wire_2129[ 11 ];
	assign fresh_wire_2132[ 12 ] = fresh_wire_2129[ 12 ];
	assign fresh_wire_2132[ 13 ] = fresh_wire_2129[ 13 ];
	assign fresh_wire_2132[ 14 ] = fresh_wire_2129[ 14 ];
	assign fresh_wire_2132[ 15 ] = fresh_wire_2129[ 15 ];
	assign fresh_wire_2132[ 16 ] = fresh_wire_2129[ 16 ];
	assign fresh_wire_2133[ 0 ] = fresh_wire_2131[ 0 ];
	assign fresh_wire_2133[ 1 ] = fresh_wire_2131[ 1 ];
	assign fresh_wire_2133[ 2 ] = fresh_wire_2131[ 2 ];
	assign fresh_wire_2133[ 3 ] = fresh_wire_2131[ 3 ];
	assign fresh_wire_2133[ 4 ] = fresh_wire_2131[ 4 ];
	assign fresh_wire_2133[ 5 ] = fresh_wire_2131[ 5 ];
	assign fresh_wire_2133[ 6 ] = fresh_wire_2131[ 6 ];
	assign fresh_wire_2133[ 7 ] = fresh_wire_2131[ 7 ];
	assign fresh_wire_2133[ 8 ] = fresh_wire_2131[ 8 ];
	assign fresh_wire_2133[ 9 ] = fresh_wire_2131[ 9 ];
	assign fresh_wire_2133[ 10 ] = fresh_wire_2131[ 10 ];
	assign fresh_wire_2133[ 11 ] = fresh_wire_2131[ 11 ];
	assign fresh_wire_2133[ 12 ] = fresh_wire_2131[ 12 ];
	assign fresh_wire_2133[ 13 ] = fresh_wire_2131[ 13 ];
	assign fresh_wire_2133[ 14 ] = fresh_wire_2131[ 14 ];
	assign fresh_wire_2133[ 15 ] = fresh_wire_2131[ 15 ];
	assign fresh_wire_2133[ 16 ] = fresh_wire_2131[ 16 ];
	assign fresh_wire_2135[ 0 ] = fresh_wire_2134[ 0 ];
	assign fresh_wire_2135[ 1 ] = fresh_wire_2134[ 1 ];
	assign fresh_wire_2135[ 2 ] = fresh_wire_2134[ 2 ];
	assign fresh_wire_2135[ 3 ] = fresh_wire_2134[ 3 ];
	assign fresh_wire_2135[ 4 ] = fresh_wire_2134[ 4 ];
	assign fresh_wire_2135[ 5 ] = fresh_wire_2134[ 5 ];
	assign fresh_wire_2135[ 6 ] = fresh_wire_2134[ 6 ];
	assign fresh_wire_2135[ 7 ] = fresh_wire_2134[ 7 ];
	assign fresh_wire_2135[ 8 ] = fresh_wire_2134[ 8 ];
	assign fresh_wire_2135[ 9 ] = fresh_wire_2134[ 9 ];
	assign fresh_wire_2135[ 10 ] = fresh_wire_2134[ 10 ];
	assign fresh_wire_2135[ 11 ] = fresh_wire_2134[ 11 ];
	assign fresh_wire_2135[ 12 ] = fresh_wire_2134[ 12 ];
	assign fresh_wire_2135[ 13 ] = fresh_wire_2134[ 13 ];
	assign fresh_wire_2135[ 14 ] = fresh_wire_2134[ 14 ];
	assign fresh_wire_2135[ 15 ] = fresh_wire_2134[ 15 ];
	assign fresh_wire_2135[ 16 ] = fresh_wire_2134[ 16 ];
	assign fresh_wire_2136[ 0 ] = fresh_wire_2280[ 0 ];
	assign fresh_wire_2136[ 1 ] = fresh_wire_2280[ 1 ];
	assign fresh_wire_2136[ 2 ] = fresh_wire_2280[ 2 ];
	assign fresh_wire_2136[ 3 ] = fresh_wire_2280[ 3 ];
	assign fresh_wire_2136[ 4 ] = fresh_wire_2280[ 4 ];
	assign fresh_wire_2136[ 5 ] = fresh_wire_2280[ 5 ];
	assign fresh_wire_2136[ 6 ] = fresh_wire_2280[ 6 ];
	assign fresh_wire_2136[ 7 ] = fresh_wire_2280[ 7 ];
	assign fresh_wire_2136[ 8 ] = fresh_wire_2280[ 8 ];
	assign fresh_wire_2136[ 9 ] = fresh_wire_2280[ 9 ];
	assign fresh_wire_2136[ 10 ] = fresh_wire_2280[ 10 ];
	assign fresh_wire_2136[ 11 ] = fresh_wire_2280[ 11 ];
	assign fresh_wire_2136[ 12 ] = fresh_wire_2280[ 12 ];
	assign fresh_wire_2136[ 13 ] = fresh_wire_2280[ 13 ];
	assign fresh_wire_2136[ 14 ] = fresh_wire_2280[ 14 ];
	assign fresh_wire_2136[ 15 ] = fresh_wire_2280[ 15 ];
	assign fresh_wire_2136[ 16 ] = fresh_wire_2280[ 16 ];
	assign fresh_wire_2138[ 0 ] = fresh_wire_1125[ 0 ];
	assign fresh_wire_2138[ 1 ] = fresh_wire_1125[ 1 ];
	assign fresh_wire_2138[ 2 ] = fresh_wire_1125[ 2 ];
	assign fresh_wire_2138[ 3 ] = fresh_wire_1125[ 3 ];
	assign fresh_wire_2138[ 4 ] = fresh_wire_1125[ 4 ];
	assign fresh_wire_2138[ 5 ] = fresh_wire_1125[ 5 ];
	assign fresh_wire_2138[ 6 ] = fresh_wire_1125[ 6 ];
	assign fresh_wire_2138[ 7 ] = fresh_wire_1125[ 7 ];
	assign fresh_wire_2138[ 8 ] = fresh_wire_1125[ 8 ];
	assign fresh_wire_2138[ 9 ] = fresh_wire_1125[ 9 ];
	assign fresh_wire_2138[ 10 ] = fresh_wire_1125[ 10 ];
	assign fresh_wire_2138[ 11 ] = fresh_wire_1125[ 11 ];
	assign fresh_wire_2138[ 12 ] = fresh_wire_1125[ 12 ];
	assign fresh_wire_2138[ 13 ] = fresh_wire_1125[ 13 ];
	assign fresh_wire_2138[ 14 ] = fresh_wire_1125[ 14 ];
	assign fresh_wire_2138[ 15 ] = fresh_wire_1125[ 15 ];
	assign fresh_wire_2138[ 16 ] = fresh_wire_2281[ 0 ];
	assign fresh_wire_2140[ 0 ] = fresh_wire_2139[ 0 ];
	assign fresh_wire_2140[ 1 ] = fresh_wire_2139[ 1 ];
	assign fresh_wire_2140[ 2 ] = fresh_wire_2139[ 2 ];
	assign fresh_wire_2140[ 3 ] = fresh_wire_2139[ 3 ];
	assign fresh_wire_2140[ 4 ] = fresh_wire_2139[ 4 ];
	assign fresh_wire_2140[ 5 ] = fresh_wire_2139[ 5 ];
	assign fresh_wire_2140[ 6 ] = fresh_wire_2139[ 6 ];
	assign fresh_wire_2140[ 7 ] = fresh_wire_2139[ 7 ];
	assign fresh_wire_2140[ 8 ] = fresh_wire_2139[ 8 ];
	assign fresh_wire_2140[ 9 ] = fresh_wire_2139[ 9 ];
	assign fresh_wire_2140[ 10 ] = fresh_wire_2139[ 10 ];
	assign fresh_wire_2140[ 11 ] = fresh_wire_2139[ 11 ];
	assign fresh_wire_2140[ 12 ] = fresh_wire_2139[ 12 ];
	assign fresh_wire_2140[ 13 ] = fresh_wire_2139[ 13 ];
	assign fresh_wire_2140[ 14 ] = fresh_wire_2139[ 14 ];
	assign fresh_wire_2140[ 15 ] = fresh_wire_2139[ 15 ];
	assign fresh_wire_2140[ 16 ] = fresh_wire_2139[ 16 ];
	assign fresh_wire_2140[ 17 ] = fresh_wire_2139[ 17 ];
	assign fresh_wire_2140[ 18 ] = fresh_wire_2139[ 18 ];
	assign fresh_wire_2140[ 19 ] = fresh_wire_2139[ 19 ];
	assign fresh_wire_2140[ 20 ] = fresh_wire_2139[ 20 ];
	assign fresh_wire_2140[ 21 ] = fresh_wire_2139[ 21 ];
	assign fresh_wire_2140[ 22 ] = fresh_wire_2139[ 22 ];
	assign fresh_wire_2140[ 23 ] = fresh_wire_2139[ 23 ];
	assign fresh_wire_2140[ 24 ] = fresh_wire_2139[ 24 ];
	assign fresh_wire_2140[ 25 ] = fresh_wire_2139[ 25 ];
	assign fresh_wire_2140[ 26 ] = fresh_wire_2139[ 26 ];
	assign fresh_wire_2140[ 27 ] = fresh_wire_2139[ 27 ];
	assign fresh_wire_2140[ 28 ] = fresh_wire_2139[ 28 ];
	assign fresh_wire_2140[ 29 ] = fresh_wire_2139[ 29 ];
	assign fresh_wire_2140[ 30 ] = fresh_wire_2139[ 30 ];
	assign fresh_wire_2140[ 31 ] = fresh_wire_2139[ 31 ];
	assign fresh_wire_2140[ 32 ] = fresh_wire_2139[ 32 ];
	assign fresh_wire_2140[ 33 ] = fresh_wire_2139[ 33 ];
	assign fresh_wire_2141[ 0 ] = fresh_wire_2282[ 0 ];
	assign fresh_wire_2141[ 1 ] = fresh_wire_2282[ 1 ];
	assign fresh_wire_2141[ 2 ] = fresh_wire_2282[ 2 ];
	assign fresh_wire_2141[ 3 ] = fresh_wire_2282[ 3 ];
	assign fresh_wire_2141[ 4 ] = fresh_wire_2282[ 4 ];
	assign fresh_wire_2141[ 5 ] = fresh_wire_2282[ 5 ];
	assign fresh_wire_2141[ 6 ] = fresh_wire_2282[ 6 ];
	assign fresh_wire_2141[ 7 ] = fresh_wire_2282[ 7 ];
	assign fresh_wire_2141[ 8 ] = fresh_wire_2282[ 8 ];
	assign fresh_wire_2141[ 9 ] = fresh_wire_2282[ 9 ];
	assign fresh_wire_2141[ 10 ] = fresh_wire_2282[ 10 ];
	assign fresh_wire_2141[ 11 ] = fresh_wire_2282[ 11 ];
	assign fresh_wire_2141[ 12 ] = fresh_wire_2282[ 12 ];
	assign fresh_wire_2141[ 13 ] = fresh_wire_2282[ 13 ];
	assign fresh_wire_2141[ 14 ] = fresh_wire_2282[ 14 ];
	assign fresh_wire_2141[ 15 ] = fresh_wire_2282[ 15 ];
	assign fresh_wire_2141[ 16 ] = fresh_wire_2282[ 16 ];
	assign fresh_wire_2141[ 17 ] = fresh_wire_2282[ 17 ];
	assign fresh_wire_2141[ 18 ] = fresh_wire_2282[ 18 ];
	assign fresh_wire_2141[ 19 ] = fresh_wire_2282[ 19 ];
	assign fresh_wire_2141[ 20 ] = fresh_wire_2282[ 20 ];
	assign fresh_wire_2141[ 21 ] = fresh_wire_2282[ 21 ];
	assign fresh_wire_2141[ 22 ] = fresh_wire_2282[ 22 ];
	assign fresh_wire_2141[ 23 ] = fresh_wire_2282[ 23 ];
	assign fresh_wire_2141[ 24 ] = fresh_wire_2282[ 24 ];
	assign fresh_wire_2141[ 25 ] = fresh_wire_2282[ 25 ];
	assign fresh_wire_2141[ 26 ] = fresh_wire_2282[ 26 ];
	assign fresh_wire_2141[ 27 ] = fresh_wire_2282[ 27 ];
	assign fresh_wire_2141[ 28 ] = fresh_wire_2282[ 28 ];
	assign fresh_wire_2141[ 29 ] = fresh_wire_2282[ 29 ];
	assign fresh_wire_2141[ 30 ] = fresh_wire_2282[ 30 ];
	assign fresh_wire_2141[ 31 ] = fresh_wire_2282[ 31 ];
	assign fresh_wire_2141[ 32 ] = fresh_wire_2282[ 32 ];
	assign fresh_wire_2141[ 33 ] = fresh_wire_2282[ 33 ];
	assign fresh_wire_2143[ 0 ] = fresh_wire_1125[ 0 ];
	assign fresh_wire_2143[ 1 ] = fresh_wire_1125[ 1 ];
	assign fresh_wire_2143[ 2 ] = fresh_wire_1125[ 2 ];
	assign fresh_wire_2143[ 3 ] = fresh_wire_1125[ 3 ];
	assign fresh_wire_2143[ 4 ] = fresh_wire_1125[ 4 ];
	assign fresh_wire_2143[ 5 ] = fresh_wire_1125[ 5 ];
	assign fresh_wire_2143[ 6 ] = fresh_wire_1125[ 6 ];
	assign fresh_wire_2143[ 7 ] = fresh_wire_1125[ 7 ];
	assign fresh_wire_2143[ 8 ] = fresh_wire_1125[ 8 ];
	assign fresh_wire_2143[ 9 ] = fresh_wire_1125[ 9 ];
	assign fresh_wire_2143[ 10 ] = fresh_wire_1125[ 10 ];
	assign fresh_wire_2143[ 11 ] = fresh_wire_1125[ 11 ];
	assign fresh_wire_2143[ 12 ] = fresh_wire_1125[ 12 ];
	assign fresh_wire_2143[ 13 ] = fresh_wire_1125[ 13 ];
	assign fresh_wire_2143[ 14 ] = fresh_wire_1125[ 14 ];
	assign fresh_wire_2143[ 15 ] = fresh_wire_1125[ 15 ];
	assign fresh_wire_2145[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_2146[ 0 ] = fresh_wire_2283[ 0 ];
	assign fresh_wire_2147[ 0 ] = fresh_wire_2144[ 0 ];
	assign fresh_wire_2147[ 1 ] = fresh_wire_2144[ 1 ];
	assign fresh_wire_2147[ 2 ] = fresh_wire_2144[ 2 ];
	assign fresh_wire_2147[ 3 ] = fresh_wire_2144[ 3 ];
	assign fresh_wire_2147[ 4 ] = fresh_wire_2144[ 4 ];
	assign fresh_wire_2147[ 5 ] = fresh_wire_2144[ 5 ];
	assign fresh_wire_2147[ 6 ] = fresh_wire_2144[ 6 ];
	assign fresh_wire_2147[ 7 ] = fresh_wire_2144[ 7 ];
	assign fresh_wire_2147[ 8 ] = fresh_wire_2144[ 8 ];
	assign fresh_wire_2147[ 9 ] = fresh_wire_2144[ 9 ];
	assign fresh_wire_2147[ 10 ] = fresh_wire_2144[ 10 ];
	assign fresh_wire_2147[ 11 ] = fresh_wire_2144[ 11 ];
	assign fresh_wire_2147[ 12 ] = fresh_wire_2144[ 12 ];
	assign fresh_wire_2147[ 13 ] = fresh_wire_2144[ 13 ];
	assign fresh_wire_2147[ 14 ] = fresh_wire_2144[ 14 ];
	assign fresh_wire_2147[ 15 ] = fresh_wire_2144[ 15 ];
	assign fresh_wire_2147[ 16 ] = fresh_wire_2284[ 0 ];
	assign fresh_wire_2149[ 0 ] = fresh_wire_2148[ 0 ];
	assign fresh_wire_2149[ 1 ] = fresh_wire_2148[ 1 ];
	assign fresh_wire_2149[ 2 ] = fresh_wire_2148[ 2 ];
	assign fresh_wire_2149[ 3 ] = fresh_wire_2148[ 3 ];
	assign fresh_wire_2149[ 4 ] = fresh_wire_2148[ 4 ];
	assign fresh_wire_2149[ 5 ] = fresh_wire_2148[ 5 ];
	assign fresh_wire_2149[ 6 ] = fresh_wire_2148[ 6 ];
	assign fresh_wire_2149[ 7 ] = fresh_wire_2148[ 7 ];
	assign fresh_wire_2149[ 8 ] = fresh_wire_2148[ 8 ];
	assign fresh_wire_2149[ 9 ] = fresh_wire_2148[ 9 ];
	assign fresh_wire_2149[ 10 ] = fresh_wire_2148[ 10 ];
	assign fresh_wire_2149[ 11 ] = fresh_wire_2148[ 11 ];
	assign fresh_wire_2149[ 12 ] = fresh_wire_2148[ 12 ];
	assign fresh_wire_2149[ 13 ] = fresh_wire_2148[ 13 ];
	assign fresh_wire_2149[ 14 ] = fresh_wire_2148[ 14 ];
	assign fresh_wire_2149[ 15 ] = fresh_wire_2148[ 15 ];
	assign fresh_wire_2149[ 16 ] = fresh_wire_2148[ 16 ];
	assign fresh_wire_2149[ 17 ] = fresh_wire_2148[ 17 ];
	assign fresh_wire_2149[ 18 ] = fresh_wire_2148[ 18 ];
	assign fresh_wire_2149[ 19 ] = fresh_wire_2148[ 19 ];
	assign fresh_wire_2149[ 20 ] = fresh_wire_2148[ 20 ];
	assign fresh_wire_2149[ 21 ] = fresh_wire_2148[ 21 ];
	assign fresh_wire_2149[ 22 ] = fresh_wire_2148[ 22 ];
	assign fresh_wire_2149[ 23 ] = fresh_wire_2148[ 23 ];
	assign fresh_wire_2149[ 24 ] = fresh_wire_2148[ 24 ];
	assign fresh_wire_2149[ 25 ] = fresh_wire_2148[ 25 ];
	assign fresh_wire_2149[ 26 ] = fresh_wire_2148[ 26 ];
	assign fresh_wire_2149[ 27 ] = fresh_wire_2148[ 27 ];
	assign fresh_wire_2149[ 28 ] = fresh_wire_2148[ 28 ];
	assign fresh_wire_2149[ 29 ] = fresh_wire_2148[ 29 ];
	assign fresh_wire_2149[ 30 ] = fresh_wire_2148[ 30 ];
	assign fresh_wire_2149[ 31 ] = fresh_wire_2148[ 31 ];
	assign fresh_wire_2149[ 32 ] = fresh_wire_2148[ 32 ];
	assign fresh_wire_2149[ 33 ] = fresh_wire_2148[ 33 ];
	assign fresh_wire_2150[ 0 ] = fresh_wire_2285[ 0 ];
	assign fresh_wire_2150[ 1 ] = fresh_wire_2285[ 1 ];
	assign fresh_wire_2150[ 2 ] = fresh_wire_2285[ 2 ];
	assign fresh_wire_2150[ 3 ] = fresh_wire_2285[ 3 ];
	assign fresh_wire_2150[ 4 ] = fresh_wire_2285[ 4 ];
	assign fresh_wire_2150[ 5 ] = fresh_wire_2285[ 5 ];
	assign fresh_wire_2150[ 6 ] = fresh_wire_2285[ 6 ];
	assign fresh_wire_2150[ 7 ] = fresh_wire_2285[ 7 ];
	assign fresh_wire_2150[ 8 ] = fresh_wire_2285[ 8 ];
	assign fresh_wire_2150[ 9 ] = fresh_wire_2285[ 9 ];
	assign fresh_wire_2150[ 10 ] = fresh_wire_2285[ 10 ];
	assign fresh_wire_2150[ 11 ] = fresh_wire_2285[ 11 ];
	assign fresh_wire_2150[ 12 ] = fresh_wire_2285[ 12 ];
	assign fresh_wire_2150[ 13 ] = fresh_wire_2285[ 13 ];
	assign fresh_wire_2150[ 14 ] = fresh_wire_2285[ 14 ];
	assign fresh_wire_2150[ 15 ] = fresh_wire_2285[ 15 ];
	assign fresh_wire_2150[ 16 ] = fresh_wire_2285[ 16 ];
	assign fresh_wire_2150[ 17 ] = fresh_wire_2285[ 17 ];
	assign fresh_wire_2150[ 18 ] = fresh_wire_2285[ 18 ];
	assign fresh_wire_2150[ 19 ] = fresh_wire_2285[ 19 ];
	assign fresh_wire_2150[ 20 ] = fresh_wire_2285[ 20 ];
	assign fresh_wire_2150[ 21 ] = fresh_wire_2285[ 21 ];
	assign fresh_wire_2150[ 22 ] = fresh_wire_2285[ 22 ];
	assign fresh_wire_2150[ 23 ] = fresh_wire_2285[ 23 ];
	assign fresh_wire_2150[ 24 ] = fresh_wire_2285[ 24 ];
	assign fresh_wire_2150[ 25 ] = fresh_wire_2285[ 25 ];
	assign fresh_wire_2150[ 26 ] = fresh_wire_2285[ 26 ];
	assign fresh_wire_2150[ 27 ] = fresh_wire_2285[ 27 ];
	assign fresh_wire_2150[ 28 ] = fresh_wire_2285[ 28 ];
	assign fresh_wire_2150[ 29 ] = fresh_wire_2285[ 29 ];
	assign fresh_wire_2150[ 30 ] = fresh_wire_2285[ 30 ];
	assign fresh_wire_2150[ 31 ] = fresh_wire_2285[ 31 ];
	assign fresh_wire_2150[ 32 ] = fresh_wire_2285[ 32 ];
	assign fresh_wire_2150[ 33 ] = fresh_wire_2285[ 33 ];
	assign fresh_wire_2152[ 0 ] = fresh_wire_2127[ 0 ];
	assign fresh_wire_2152[ 1 ] = fresh_wire_2127[ 1 ];
	assign fresh_wire_2152[ 2 ] = fresh_wire_2127[ 2 ];
	assign fresh_wire_2152[ 3 ] = fresh_wire_2127[ 3 ];
	assign fresh_wire_2152[ 4 ] = fresh_wire_2127[ 4 ];
	assign fresh_wire_2152[ 5 ] = fresh_wire_2127[ 5 ];
	assign fresh_wire_2152[ 6 ] = fresh_wire_2127[ 6 ];
	assign fresh_wire_2152[ 7 ] = fresh_wire_2127[ 7 ];
	assign fresh_wire_2152[ 8 ] = fresh_wire_2127[ 8 ];
	assign fresh_wire_2152[ 9 ] = fresh_wire_2127[ 9 ];
	assign fresh_wire_2152[ 10 ] = fresh_wire_2127[ 10 ];
	assign fresh_wire_2152[ 11 ] = fresh_wire_2127[ 11 ];
	assign fresh_wire_2152[ 12 ] = fresh_wire_2127[ 12 ];
	assign fresh_wire_2152[ 13 ] = fresh_wire_2127[ 13 ];
	assign fresh_wire_2152[ 14 ] = fresh_wire_2127[ 14 ];
	assign fresh_wire_2152[ 15 ] = fresh_wire_2127[ 15 ];
	assign fresh_wire_2154[ 0 ] = fresh_wire_2116[ 0 ];
	assign fresh_wire_2154[ 1 ] = fresh_wire_2116[ 1 ];
	assign fresh_wire_2154[ 2 ] = fresh_wire_2116[ 2 ];
	assign fresh_wire_2154[ 3 ] = fresh_wire_2116[ 3 ];
	assign fresh_wire_2154[ 4 ] = fresh_wire_2116[ 4 ];
	assign fresh_wire_2154[ 5 ] = fresh_wire_2116[ 5 ];
	assign fresh_wire_2154[ 6 ] = fresh_wire_2116[ 6 ];
	assign fresh_wire_2154[ 7 ] = fresh_wire_2116[ 7 ];
	assign fresh_wire_2154[ 8 ] = fresh_wire_2116[ 8 ];
	assign fresh_wire_2154[ 9 ] = fresh_wire_2116[ 9 ];
	assign fresh_wire_2154[ 10 ] = fresh_wire_2116[ 10 ];
	assign fresh_wire_2154[ 11 ] = fresh_wire_2116[ 11 ];
	assign fresh_wire_2154[ 12 ] = fresh_wire_2116[ 12 ];
	assign fresh_wire_2154[ 13 ] = fresh_wire_2116[ 13 ];
	assign fresh_wire_2154[ 14 ] = fresh_wire_2116[ 14 ];
	assign fresh_wire_2154[ 15 ] = fresh_wire_2116[ 15 ];
	assign fresh_wire_2156[ 0 ] = fresh_wire_2153[ 0 ];
	assign fresh_wire_2156[ 1 ] = fresh_wire_2153[ 1 ];
	assign fresh_wire_2156[ 2 ] = fresh_wire_2153[ 2 ];
	assign fresh_wire_2156[ 3 ] = fresh_wire_2153[ 3 ];
	assign fresh_wire_2156[ 4 ] = fresh_wire_2153[ 4 ];
	assign fresh_wire_2156[ 5 ] = fresh_wire_2153[ 5 ];
	assign fresh_wire_2156[ 6 ] = fresh_wire_2153[ 6 ];
	assign fresh_wire_2156[ 7 ] = fresh_wire_2153[ 7 ];
	assign fresh_wire_2156[ 8 ] = fresh_wire_2153[ 8 ];
	assign fresh_wire_2156[ 9 ] = fresh_wire_2153[ 9 ];
	assign fresh_wire_2156[ 10 ] = fresh_wire_2153[ 10 ];
	assign fresh_wire_2156[ 11 ] = fresh_wire_2153[ 11 ];
	assign fresh_wire_2156[ 12 ] = fresh_wire_2153[ 12 ];
	assign fresh_wire_2156[ 13 ] = fresh_wire_2153[ 13 ];
	assign fresh_wire_2156[ 14 ] = fresh_wire_2153[ 14 ];
	assign fresh_wire_2156[ 15 ] = fresh_wire_2153[ 15 ];
	assign fresh_wire_2156[ 16 ] = fresh_wire_2153[ 16 ];
	assign fresh_wire_2157[ 0 ] = fresh_wire_2155[ 0 ];
	assign fresh_wire_2157[ 1 ] = fresh_wire_2155[ 1 ];
	assign fresh_wire_2157[ 2 ] = fresh_wire_2155[ 2 ];
	assign fresh_wire_2157[ 3 ] = fresh_wire_2155[ 3 ];
	assign fresh_wire_2157[ 4 ] = fresh_wire_2155[ 4 ];
	assign fresh_wire_2157[ 5 ] = fresh_wire_2155[ 5 ];
	assign fresh_wire_2157[ 6 ] = fresh_wire_2155[ 6 ];
	assign fresh_wire_2157[ 7 ] = fresh_wire_2155[ 7 ];
	assign fresh_wire_2157[ 8 ] = fresh_wire_2155[ 8 ];
	assign fresh_wire_2157[ 9 ] = fresh_wire_2155[ 9 ];
	assign fresh_wire_2157[ 10 ] = fresh_wire_2155[ 10 ];
	assign fresh_wire_2157[ 11 ] = fresh_wire_2155[ 11 ];
	assign fresh_wire_2157[ 12 ] = fresh_wire_2155[ 12 ];
	assign fresh_wire_2157[ 13 ] = fresh_wire_2155[ 13 ];
	assign fresh_wire_2157[ 14 ] = fresh_wire_2155[ 14 ];
	assign fresh_wire_2157[ 15 ] = fresh_wire_2155[ 15 ];
	assign fresh_wire_2157[ 16 ] = fresh_wire_2155[ 16 ];
	assign fresh_wire_2159[ 0 ] = fresh_wire_2158[ 0 ];
	assign fresh_wire_2159[ 1 ] = fresh_wire_2158[ 1 ];
	assign fresh_wire_2159[ 2 ] = fresh_wire_2158[ 2 ];
	assign fresh_wire_2159[ 3 ] = fresh_wire_2158[ 3 ];
	assign fresh_wire_2159[ 4 ] = fresh_wire_2158[ 4 ];
	assign fresh_wire_2159[ 5 ] = fresh_wire_2158[ 5 ];
	assign fresh_wire_2159[ 6 ] = fresh_wire_2158[ 6 ];
	assign fresh_wire_2159[ 7 ] = fresh_wire_2158[ 7 ];
	assign fresh_wire_2159[ 8 ] = fresh_wire_2158[ 8 ];
	assign fresh_wire_2159[ 9 ] = fresh_wire_2158[ 9 ];
	assign fresh_wire_2159[ 10 ] = fresh_wire_2158[ 10 ];
	assign fresh_wire_2159[ 11 ] = fresh_wire_2158[ 11 ];
	assign fresh_wire_2159[ 12 ] = fresh_wire_2158[ 12 ];
	assign fresh_wire_2159[ 13 ] = fresh_wire_2158[ 13 ];
	assign fresh_wire_2159[ 14 ] = fresh_wire_2158[ 14 ];
	assign fresh_wire_2159[ 15 ] = fresh_wire_2158[ 15 ];
	assign fresh_wire_2159[ 16 ] = fresh_wire_2158[ 16 ];
	assign fresh_wire_2160[ 0 ] = fresh_wire_2286[ 0 ];
	assign fresh_wire_2160[ 1 ] = fresh_wire_2286[ 1 ];
	assign fresh_wire_2160[ 2 ] = fresh_wire_2286[ 2 ];
	assign fresh_wire_2160[ 3 ] = fresh_wire_2286[ 3 ];
	assign fresh_wire_2160[ 4 ] = fresh_wire_2286[ 4 ];
	assign fresh_wire_2160[ 5 ] = fresh_wire_2286[ 5 ];
	assign fresh_wire_2160[ 6 ] = fresh_wire_2286[ 6 ];
	assign fresh_wire_2160[ 7 ] = fresh_wire_2286[ 7 ];
	assign fresh_wire_2160[ 8 ] = fresh_wire_2286[ 8 ];
	assign fresh_wire_2160[ 9 ] = fresh_wire_2286[ 9 ];
	assign fresh_wire_2160[ 10 ] = fresh_wire_2286[ 10 ];
	assign fresh_wire_2160[ 11 ] = fresh_wire_2286[ 11 ];
	assign fresh_wire_2160[ 12 ] = fresh_wire_2286[ 12 ];
	assign fresh_wire_2160[ 13 ] = fresh_wire_2286[ 13 ];
	assign fresh_wire_2160[ 14 ] = fresh_wire_2286[ 14 ];
	assign fresh_wire_2160[ 15 ] = fresh_wire_2286[ 15 ];
	assign fresh_wire_2160[ 16 ] = fresh_wire_2286[ 16 ];
	assign fresh_wire_2162[ 0 ] = fresh_wire_2176[ 0 ];
	assign fresh_wire_2162[ 1 ] = fresh_wire_2176[ 1 ];
	assign fresh_wire_2162[ 2 ] = fresh_wire_2176[ 2 ];
	assign fresh_wire_2162[ 3 ] = fresh_wire_2176[ 3 ];
	assign fresh_wire_2162[ 4 ] = fresh_wire_2176[ 4 ];
	assign fresh_wire_2162[ 5 ] = fresh_wire_2176[ 5 ];
	assign fresh_wire_2162[ 6 ] = fresh_wire_2176[ 6 ];
	assign fresh_wire_2162[ 7 ] = fresh_wire_2176[ 7 ];
	assign fresh_wire_2162[ 8 ] = fresh_wire_2176[ 8 ];
	assign fresh_wire_2162[ 9 ] = fresh_wire_2176[ 9 ];
	assign fresh_wire_2162[ 10 ] = fresh_wire_2176[ 10 ];
	assign fresh_wire_2162[ 11 ] = fresh_wire_2176[ 11 ];
	assign fresh_wire_2162[ 12 ] = fresh_wire_2176[ 12 ];
	assign fresh_wire_2162[ 13 ] = fresh_wire_2176[ 13 ];
	assign fresh_wire_2162[ 14 ] = fresh_wire_2176[ 14 ];
	assign fresh_wire_2162[ 15 ] = fresh_wire_2176[ 15 ];
	assign fresh_wire_2164[ 0 ] = fresh_wire_2248[ 0 ];
	assign fresh_wire_2164[ 1 ] = fresh_wire_2248[ 1 ];
	assign fresh_wire_2164[ 2 ] = fresh_wire_2248[ 2 ];
	assign fresh_wire_2164[ 3 ] = fresh_wire_2248[ 3 ];
	assign fresh_wire_2164[ 4 ] = fresh_wire_2248[ 4 ];
	assign fresh_wire_2164[ 5 ] = fresh_wire_2248[ 5 ];
	assign fresh_wire_2164[ 6 ] = fresh_wire_2248[ 6 ];
	assign fresh_wire_2164[ 7 ] = fresh_wire_2248[ 7 ];
	assign fresh_wire_2164[ 8 ] = fresh_wire_2248[ 8 ];
	assign fresh_wire_2164[ 9 ] = fresh_wire_2248[ 9 ];
	assign fresh_wire_2164[ 10 ] = fresh_wire_2248[ 10 ];
	assign fresh_wire_2164[ 11 ] = fresh_wire_2248[ 11 ];
	assign fresh_wire_2164[ 12 ] = fresh_wire_2248[ 12 ];
	assign fresh_wire_2164[ 13 ] = fresh_wire_2248[ 13 ];
	assign fresh_wire_2164[ 14 ] = fresh_wire_2248[ 14 ];
	assign fresh_wire_2164[ 15 ] = fresh_wire_2248[ 15 ];
	assign fresh_wire_2166[ 0 ] = fresh_wire_2163[ 0 ];
	assign fresh_wire_2166[ 1 ] = fresh_wire_2163[ 1 ];
	assign fresh_wire_2166[ 2 ] = fresh_wire_2163[ 2 ];
	assign fresh_wire_2166[ 3 ] = fresh_wire_2163[ 3 ];
	assign fresh_wire_2166[ 4 ] = fresh_wire_2163[ 4 ];
	assign fresh_wire_2166[ 5 ] = fresh_wire_2163[ 5 ];
	assign fresh_wire_2166[ 6 ] = fresh_wire_2163[ 6 ];
	assign fresh_wire_2166[ 7 ] = fresh_wire_2163[ 7 ];
	assign fresh_wire_2166[ 8 ] = fresh_wire_2163[ 8 ];
	assign fresh_wire_2166[ 9 ] = fresh_wire_2163[ 9 ];
	assign fresh_wire_2166[ 10 ] = fresh_wire_2163[ 10 ];
	assign fresh_wire_2166[ 11 ] = fresh_wire_2163[ 11 ];
	assign fresh_wire_2166[ 12 ] = fresh_wire_2163[ 12 ];
	assign fresh_wire_2166[ 13 ] = fresh_wire_2163[ 13 ];
	assign fresh_wire_2166[ 14 ] = fresh_wire_2163[ 14 ];
	assign fresh_wire_2166[ 15 ] = fresh_wire_2163[ 15 ];
	assign fresh_wire_2166[ 16 ] = fresh_wire_2163[ 16 ];
	assign fresh_wire_2167[ 0 ] = fresh_wire_2165[ 0 ];
	assign fresh_wire_2167[ 1 ] = fresh_wire_2165[ 1 ];
	assign fresh_wire_2167[ 2 ] = fresh_wire_2165[ 2 ];
	assign fresh_wire_2167[ 3 ] = fresh_wire_2165[ 3 ];
	assign fresh_wire_2167[ 4 ] = fresh_wire_2165[ 4 ];
	assign fresh_wire_2167[ 5 ] = fresh_wire_2165[ 5 ];
	assign fresh_wire_2167[ 6 ] = fresh_wire_2165[ 6 ];
	assign fresh_wire_2167[ 7 ] = fresh_wire_2165[ 7 ];
	assign fresh_wire_2167[ 8 ] = fresh_wire_2165[ 8 ];
	assign fresh_wire_2167[ 9 ] = fresh_wire_2165[ 9 ];
	assign fresh_wire_2167[ 10 ] = fresh_wire_2165[ 10 ];
	assign fresh_wire_2167[ 11 ] = fresh_wire_2165[ 11 ];
	assign fresh_wire_2167[ 12 ] = fresh_wire_2165[ 12 ];
	assign fresh_wire_2167[ 13 ] = fresh_wire_2165[ 13 ];
	assign fresh_wire_2167[ 14 ] = fresh_wire_2165[ 14 ];
	assign fresh_wire_2167[ 15 ] = fresh_wire_2165[ 15 ];
	assign fresh_wire_2167[ 16 ] = fresh_wire_2165[ 16 ];
	assign fresh_wire_2169[ 0 ] = fresh_wire_2168[ 0 ];
	assign fresh_wire_2169[ 1 ] = fresh_wire_2168[ 1 ];
	assign fresh_wire_2169[ 2 ] = fresh_wire_2168[ 2 ];
	assign fresh_wire_2169[ 3 ] = fresh_wire_2168[ 3 ];
	assign fresh_wire_2169[ 4 ] = fresh_wire_2168[ 4 ];
	assign fresh_wire_2169[ 5 ] = fresh_wire_2168[ 5 ];
	assign fresh_wire_2169[ 6 ] = fresh_wire_2168[ 6 ];
	assign fresh_wire_2169[ 7 ] = fresh_wire_2168[ 7 ];
	assign fresh_wire_2169[ 8 ] = fresh_wire_2168[ 8 ];
	assign fresh_wire_2169[ 9 ] = fresh_wire_2168[ 9 ];
	assign fresh_wire_2169[ 10 ] = fresh_wire_2168[ 10 ];
	assign fresh_wire_2169[ 11 ] = fresh_wire_2168[ 11 ];
	assign fresh_wire_2169[ 12 ] = fresh_wire_2168[ 12 ];
	assign fresh_wire_2169[ 13 ] = fresh_wire_2168[ 13 ];
	assign fresh_wire_2169[ 14 ] = fresh_wire_2168[ 14 ];
	assign fresh_wire_2169[ 15 ] = fresh_wire_2168[ 15 ];
	assign fresh_wire_2169[ 16 ] = fresh_wire_2168[ 16 ];
	assign fresh_wire_2170[ 0 ] = fresh_wire_2287[ 0 ];
	assign fresh_wire_2170[ 1 ] = fresh_wire_2287[ 1 ];
	assign fresh_wire_2170[ 2 ] = fresh_wire_2287[ 2 ];
	assign fresh_wire_2170[ 3 ] = fresh_wire_2287[ 3 ];
	assign fresh_wire_2170[ 4 ] = fresh_wire_2287[ 4 ];
	assign fresh_wire_2170[ 5 ] = fresh_wire_2287[ 5 ];
	assign fresh_wire_2170[ 6 ] = fresh_wire_2287[ 6 ];
	assign fresh_wire_2170[ 7 ] = fresh_wire_2287[ 7 ];
	assign fresh_wire_2170[ 8 ] = fresh_wire_2287[ 8 ];
	assign fresh_wire_2170[ 9 ] = fresh_wire_2287[ 9 ];
	assign fresh_wire_2170[ 10 ] = fresh_wire_2287[ 10 ];
	assign fresh_wire_2170[ 11 ] = fresh_wire_2287[ 11 ];
	assign fresh_wire_2170[ 12 ] = fresh_wire_2287[ 12 ];
	assign fresh_wire_2170[ 13 ] = fresh_wire_2287[ 13 ];
	assign fresh_wire_2170[ 14 ] = fresh_wire_2287[ 14 ];
	assign fresh_wire_2170[ 15 ] = fresh_wire_2287[ 15 ];
	assign fresh_wire_2170[ 16 ] = fresh_wire_2287[ 16 ];
	assign fresh_wire_2172[ 0 ] = fresh_wire_1581[ 0 ];
	assign fresh_wire_2172[ 1 ] = fresh_wire_1581[ 1 ];
	assign fresh_wire_2172[ 2 ] = fresh_wire_1581[ 2 ];
	assign fresh_wire_2172[ 3 ] = fresh_wire_1581[ 3 ];
	assign fresh_wire_2172[ 4 ] = fresh_wire_1581[ 4 ];
	assign fresh_wire_2172[ 5 ] = fresh_wire_1581[ 5 ];
	assign fresh_wire_2172[ 6 ] = fresh_wire_1581[ 6 ];
	assign fresh_wire_2172[ 7 ] = fresh_wire_1581[ 7 ];
	assign fresh_wire_2172[ 8 ] = fresh_wire_1581[ 8 ];
	assign fresh_wire_2172[ 9 ] = fresh_wire_1581[ 9 ];
	assign fresh_wire_2172[ 10 ] = fresh_wire_1581[ 10 ];
	assign fresh_wire_2172[ 11 ] = fresh_wire_1581[ 11 ];
	assign fresh_wire_2172[ 12 ] = fresh_wire_1581[ 12 ];
	assign fresh_wire_2172[ 13 ] = fresh_wire_1581[ 13 ];
	assign fresh_wire_2172[ 14 ] = fresh_wire_1581[ 14 ];
	assign fresh_wire_2172[ 15 ] = fresh_wire_1581[ 15 ];
	assign fresh_wire_2172[ 16 ] = fresh_wire_2288[ 0 ];
	assign fresh_wire_2174[ 0 ] = fresh_wire_2173[ 0 ];
	assign fresh_wire_2174[ 1 ] = fresh_wire_2173[ 1 ];
	assign fresh_wire_2174[ 2 ] = fresh_wire_2173[ 2 ];
	assign fresh_wire_2174[ 3 ] = fresh_wire_2173[ 3 ];
	assign fresh_wire_2174[ 4 ] = fresh_wire_2173[ 4 ];
	assign fresh_wire_2174[ 5 ] = fresh_wire_2173[ 5 ];
	assign fresh_wire_2174[ 6 ] = fresh_wire_2173[ 6 ];
	assign fresh_wire_2174[ 7 ] = fresh_wire_2173[ 7 ];
	assign fresh_wire_2174[ 8 ] = fresh_wire_2173[ 8 ];
	assign fresh_wire_2174[ 9 ] = fresh_wire_2173[ 9 ];
	assign fresh_wire_2174[ 10 ] = fresh_wire_2173[ 10 ];
	assign fresh_wire_2174[ 11 ] = fresh_wire_2173[ 11 ];
	assign fresh_wire_2174[ 12 ] = fresh_wire_2173[ 12 ];
	assign fresh_wire_2174[ 13 ] = fresh_wire_2173[ 13 ];
	assign fresh_wire_2174[ 14 ] = fresh_wire_2173[ 14 ];
	assign fresh_wire_2174[ 15 ] = fresh_wire_2173[ 15 ];
	assign fresh_wire_2174[ 16 ] = fresh_wire_2173[ 16 ];
	assign fresh_wire_2174[ 17 ] = fresh_wire_2173[ 17 ];
	assign fresh_wire_2174[ 18 ] = fresh_wire_2173[ 18 ];
	assign fresh_wire_2174[ 19 ] = fresh_wire_2173[ 19 ];
	assign fresh_wire_2174[ 20 ] = fresh_wire_2173[ 20 ];
	assign fresh_wire_2174[ 21 ] = fresh_wire_2173[ 21 ];
	assign fresh_wire_2174[ 22 ] = fresh_wire_2173[ 22 ];
	assign fresh_wire_2174[ 23 ] = fresh_wire_2173[ 23 ];
	assign fresh_wire_2174[ 24 ] = fresh_wire_2173[ 24 ];
	assign fresh_wire_2174[ 25 ] = fresh_wire_2173[ 25 ];
	assign fresh_wire_2174[ 26 ] = fresh_wire_2173[ 26 ];
	assign fresh_wire_2174[ 27 ] = fresh_wire_2173[ 27 ];
	assign fresh_wire_2174[ 28 ] = fresh_wire_2173[ 28 ];
	assign fresh_wire_2174[ 29 ] = fresh_wire_2173[ 29 ];
	assign fresh_wire_2174[ 30 ] = fresh_wire_2173[ 30 ];
	assign fresh_wire_2174[ 31 ] = fresh_wire_2173[ 31 ];
	assign fresh_wire_2174[ 32 ] = fresh_wire_2173[ 32 ];
	assign fresh_wire_2174[ 33 ] = fresh_wire_2173[ 33 ];
	assign fresh_wire_2175[ 0 ] = fresh_wire_2289[ 0 ];
	assign fresh_wire_2175[ 1 ] = fresh_wire_2289[ 1 ];
	assign fresh_wire_2175[ 2 ] = fresh_wire_2289[ 2 ];
	assign fresh_wire_2175[ 3 ] = fresh_wire_2289[ 3 ];
	assign fresh_wire_2175[ 4 ] = fresh_wire_2289[ 4 ];
	assign fresh_wire_2175[ 5 ] = fresh_wire_2289[ 5 ];
	assign fresh_wire_2175[ 6 ] = fresh_wire_2289[ 6 ];
	assign fresh_wire_2175[ 7 ] = fresh_wire_2289[ 7 ];
	assign fresh_wire_2175[ 8 ] = fresh_wire_2289[ 8 ];
	assign fresh_wire_2175[ 9 ] = fresh_wire_2289[ 9 ];
	assign fresh_wire_2175[ 10 ] = fresh_wire_2289[ 10 ];
	assign fresh_wire_2175[ 11 ] = fresh_wire_2289[ 11 ];
	assign fresh_wire_2175[ 12 ] = fresh_wire_2289[ 12 ];
	assign fresh_wire_2175[ 13 ] = fresh_wire_2289[ 13 ];
	assign fresh_wire_2175[ 14 ] = fresh_wire_2289[ 14 ];
	assign fresh_wire_2175[ 15 ] = fresh_wire_2289[ 15 ];
	assign fresh_wire_2175[ 16 ] = fresh_wire_2289[ 16 ];
	assign fresh_wire_2175[ 17 ] = fresh_wire_2289[ 17 ];
	assign fresh_wire_2175[ 18 ] = fresh_wire_2289[ 18 ];
	assign fresh_wire_2175[ 19 ] = fresh_wire_2289[ 19 ];
	assign fresh_wire_2175[ 20 ] = fresh_wire_2289[ 20 ];
	assign fresh_wire_2175[ 21 ] = fresh_wire_2289[ 21 ];
	assign fresh_wire_2175[ 22 ] = fresh_wire_2289[ 22 ];
	assign fresh_wire_2175[ 23 ] = fresh_wire_2289[ 23 ];
	assign fresh_wire_2175[ 24 ] = fresh_wire_2289[ 24 ];
	assign fresh_wire_2175[ 25 ] = fresh_wire_2289[ 25 ];
	assign fresh_wire_2175[ 26 ] = fresh_wire_2289[ 26 ];
	assign fresh_wire_2175[ 27 ] = fresh_wire_2289[ 27 ];
	assign fresh_wire_2175[ 28 ] = fresh_wire_2289[ 28 ];
	assign fresh_wire_2175[ 29 ] = fresh_wire_2289[ 29 ];
	assign fresh_wire_2175[ 30 ] = fresh_wire_2289[ 30 ];
	assign fresh_wire_2175[ 31 ] = fresh_wire_2289[ 31 ];
	assign fresh_wire_2175[ 32 ] = fresh_wire_2289[ 32 ];
	assign fresh_wire_2175[ 33 ] = fresh_wire_2289[ 33 ];
	assign fresh_wire_2178[ 0 ] = fresh_wire_2229[ 0 ];
	assign fresh_wire_2178[ 1 ] = fresh_wire_2229[ 1 ];
	assign fresh_wire_2178[ 2 ] = fresh_wire_2229[ 2 ];
	assign fresh_wire_2178[ 3 ] = fresh_wire_2229[ 3 ];
	assign fresh_wire_2178[ 4 ] = fresh_wire_2229[ 4 ];
	assign fresh_wire_2178[ 5 ] = fresh_wire_2229[ 5 ];
	assign fresh_wire_2178[ 6 ] = fresh_wire_2229[ 6 ];
	assign fresh_wire_2178[ 7 ] = fresh_wire_2229[ 7 ];
	assign fresh_wire_2178[ 8 ] = fresh_wire_2229[ 8 ];
	assign fresh_wire_2178[ 9 ] = fresh_wire_2229[ 9 ];
	assign fresh_wire_2178[ 10 ] = fresh_wire_2229[ 10 ];
	assign fresh_wire_2178[ 11 ] = fresh_wire_2229[ 11 ];
	assign fresh_wire_2178[ 12 ] = fresh_wire_2229[ 12 ];
	assign fresh_wire_2178[ 13 ] = fresh_wire_2229[ 13 ];
	assign fresh_wire_2178[ 14 ] = fresh_wire_2229[ 14 ];
	assign fresh_wire_2178[ 15 ] = fresh_wire_2229[ 15 ];
	assign fresh_wire_2180[ 0 ] = fresh_wire_2179[ 0 ];
	assign fresh_wire_2180[ 1 ] = fresh_wire_2179[ 1 ];
	assign fresh_wire_2180[ 2 ] = fresh_wire_2179[ 2 ];
	assign fresh_wire_2180[ 3 ] = fresh_wire_2179[ 3 ];
	assign fresh_wire_2180[ 4 ] = fresh_wire_2179[ 4 ];
	assign fresh_wire_2180[ 5 ] = fresh_wire_2179[ 5 ];
	assign fresh_wire_2180[ 6 ] = fresh_wire_2179[ 6 ];
	assign fresh_wire_2180[ 7 ] = fresh_wire_2179[ 7 ];
	assign fresh_wire_2180[ 8 ] = fresh_wire_2179[ 8 ];
	assign fresh_wire_2180[ 9 ] = fresh_wire_2179[ 9 ];
	assign fresh_wire_2180[ 10 ] = fresh_wire_2179[ 10 ];
	assign fresh_wire_2180[ 11 ] = fresh_wire_2179[ 11 ];
	assign fresh_wire_2180[ 12 ] = fresh_wire_2179[ 12 ];
	assign fresh_wire_2180[ 13 ] = fresh_wire_2179[ 13 ];
	assign fresh_wire_2180[ 14 ] = fresh_wire_2179[ 14 ];
	assign fresh_wire_2180[ 15 ] = fresh_wire_2179[ 15 ];
	assign fresh_wire_2180[ 16 ] = fresh_wire_2179[ 16 ];
	assign fresh_wire_2181[ 0 ] = fresh_wire_2295[ 0 ];
	assign fresh_wire_2181[ 1 ] = fresh_wire_2295[ 1 ];
	assign fresh_wire_2181[ 2 ] = fresh_wire_2295[ 2 ];
	assign fresh_wire_2181[ 3 ] = fresh_wire_2295[ 3 ];
	assign fresh_wire_2181[ 4 ] = fresh_wire_2295[ 4 ];
	assign fresh_wire_2181[ 5 ] = fresh_wire_2295[ 5 ];
	assign fresh_wire_2181[ 6 ] = fresh_wire_2295[ 6 ];
	assign fresh_wire_2181[ 7 ] = fresh_wire_2295[ 7 ];
	assign fresh_wire_2181[ 8 ] = fresh_wire_2295[ 8 ];
	assign fresh_wire_2181[ 9 ] = fresh_wire_2295[ 9 ];
	assign fresh_wire_2181[ 10 ] = fresh_wire_2295[ 10 ];
	assign fresh_wire_2181[ 11 ] = fresh_wire_2295[ 11 ];
	assign fresh_wire_2181[ 12 ] = fresh_wire_2295[ 12 ];
	assign fresh_wire_2181[ 13 ] = fresh_wire_2295[ 13 ];
	assign fresh_wire_2181[ 14 ] = fresh_wire_2295[ 14 ];
	assign fresh_wire_2181[ 15 ] = fresh_wire_2295[ 15 ];
	assign fresh_wire_2181[ 16 ] = fresh_wire_2295[ 16 ];
	assign fresh_wire_2183[ 0 ] = fresh_wire_2182[ 0 ];
	assign fresh_wire_2183[ 1 ] = fresh_wire_2182[ 1 ];
	assign fresh_wire_2183[ 2 ] = fresh_wire_2182[ 2 ];
	assign fresh_wire_2183[ 3 ] = fresh_wire_2182[ 3 ];
	assign fresh_wire_2183[ 4 ] = fresh_wire_2182[ 4 ];
	assign fresh_wire_2183[ 5 ] = fresh_wire_2182[ 5 ];
	assign fresh_wire_2183[ 6 ] = fresh_wire_2182[ 6 ];
	assign fresh_wire_2183[ 7 ] = fresh_wire_2182[ 7 ];
	assign fresh_wire_2183[ 8 ] = fresh_wire_2182[ 8 ];
	assign fresh_wire_2183[ 9 ] = fresh_wire_2182[ 9 ];
	assign fresh_wire_2183[ 10 ] = fresh_wire_2182[ 10 ];
	assign fresh_wire_2183[ 11 ] = fresh_wire_2182[ 11 ];
	assign fresh_wire_2183[ 12 ] = fresh_wire_2182[ 12 ];
	assign fresh_wire_2183[ 13 ] = fresh_wire_2182[ 13 ];
	assign fresh_wire_2183[ 14 ] = fresh_wire_2182[ 14 ];
	assign fresh_wire_2183[ 15 ] = fresh_wire_2182[ 15 ];
	assign fresh_wire_2183[ 16 ] = fresh_wire_2182[ 16 ];
	assign fresh_wire_2184[ 0 ] = fresh_wire_2294[ 0 ];
	assign fresh_wire_2184[ 1 ] = fresh_wire_2294[ 1 ];
	assign fresh_wire_2184[ 2 ] = fresh_wire_2294[ 2 ];
	assign fresh_wire_2184[ 3 ] = fresh_wire_2294[ 3 ];
	assign fresh_wire_2184[ 4 ] = fresh_wire_2294[ 4 ];
	assign fresh_wire_2184[ 5 ] = fresh_wire_2294[ 5 ];
	assign fresh_wire_2184[ 6 ] = fresh_wire_2294[ 6 ];
	assign fresh_wire_2184[ 7 ] = fresh_wire_2294[ 7 ];
	assign fresh_wire_2184[ 8 ] = fresh_wire_2294[ 8 ];
	assign fresh_wire_2184[ 9 ] = fresh_wire_2294[ 9 ];
	assign fresh_wire_2184[ 10 ] = fresh_wire_2294[ 10 ];
	assign fresh_wire_2184[ 11 ] = fresh_wire_2294[ 11 ];
	assign fresh_wire_2184[ 12 ] = fresh_wire_2294[ 12 ];
	assign fresh_wire_2184[ 13 ] = fresh_wire_2294[ 13 ];
	assign fresh_wire_2184[ 14 ] = fresh_wire_2294[ 14 ];
	assign fresh_wire_2184[ 15 ] = fresh_wire_2294[ 15 ];
	assign fresh_wire_2184[ 16 ] = fresh_wire_2294[ 16 ];
	assign fresh_wire_2186[ 0 ] = fresh_wire_2161[ 0 ];
	assign fresh_wire_2186[ 1 ] = fresh_wire_2161[ 1 ];
	assign fresh_wire_2186[ 2 ] = fresh_wire_2161[ 2 ];
	assign fresh_wire_2186[ 3 ] = fresh_wire_2161[ 3 ];
	assign fresh_wire_2186[ 4 ] = fresh_wire_2161[ 4 ];
	assign fresh_wire_2186[ 5 ] = fresh_wire_2161[ 5 ];
	assign fresh_wire_2186[ 6 ] = fresh_wire_2161[ 6 ];
	assign fresh_wire_2186[ 7 ] = fresh_wire_2161[ 7 ];
	assign fresh_wire_2186[ 8 ] = fresh_wire_2161[ 8 ];
	assign fresh_wire_2186[ 9 ] = fresh_wire_2161[ 9 ];
	assign fresh_wire_2186[ 10 ] = fresh_wire_2161[ 10 ];
	assign fresh_wire_2186[ 11 ] = fresh_wire_2161[ 11 ];
	assign fresh_wire_2186[ 12 ] = fresh_wire_2161[ 12 ];
	assign fresh_wire_2186[ 13 ] = fresh_wire_2161[ 13 ];
	assign fresh_wire_2186[ 14 ] = fresh_wire_2161[ 14 ];
	assign fresh_wire_2186[ 15 ] = fresh_wire_2161[ 15 ];
	assign fresh_wire_2188[ 0 ] = fresh_wire_2238[ 0 ];
	assign fresh_wire_2188[ 1 ] = fresh_wire_2238[ 1 ];
	assign fresh_wire_2188[ 2 ] = fresh_wire_2238[ 2 ];
	assign fresh_wire_2188[ 3 ] = fresh_wire_2238[ 3 ];
	assign fresh_wire_2188[ 4 ] = fresh_wire_2238[ 4 ];
	assign fresh_wire_2188[ 5 ] = fresh_wire_2238[ 5 ];
	assign fresh_wire_2188[ 6 ] = fresh_wire_2238[ 6 ];
	assign fresh_wire_2188[ 7 ] = fresh_wire_2238[ 7 ];
	assign fresh_wire_2188[ 8 ] = fresh_wire_2238[ 8 ];
	assign fresh_wire_2188[ 9 ] = fresh_wire_2238[ 9 ];
	assign fresh_wire_2188[ 10 ] = fresh_wire_2238[ 10 ];
	assign fresh_wire_2188[ 11 ] = fresh_wire_2238[ 11 ];
	assign fresh_wire_2188[ 12 ] = fresh_wire_2238[ 12 ];
	assign fresh_wire_2188[ 13 ] = fresh_wire_2238[ 13 ];
	assign fresh_wire_2188[ 14 ] = fresh_wire_2238[ 14 ];
	assign fresh_wire_2188[ 15 ] = fresh_wire_2238[ 15 ];
	assign fresh_wire_2190[ 0 ] = fresh_wire_2187[ 0 ];
	assign fresh_wire_2190[ 1 ] = fresh_wire_2187[ 1 ];
	assign fresh_wire_2190[ 2 ] = fresh_wire_2187[ 2 ];
	assign fresh_wire_2190[ 3 ] = fresh_wire_2187[ 3 ];
	assign fresh_wire_2190[ 4 ] = fresh_wire_2187[ 4 ];
	assign fresh_wire_2190[ 5 ] = fresh_wire_2187[ 5 ];
	assign fresh_wire_2190[ 6 ] = fresh_wire_2187[ 6 ];
	assign fresh_wire_2190[ 7 ] = fresh_wire_2187[ 7 ];
	assign fresh_wire_2190[ 8 ] = fresh_wire_2187[ 8 ];
	assign fresh_wire_2190[ 9 ] = fresh_wire_2187[ 9 ];
	assign fresh_wire_2190[ 10 ] = fresh_wire_2187[ 10 ];
	assign fresh_wire_2190[ 11 ] = fresh_wire_2187[ 11 ];
	assign fresh_wire_2190[ 12 ] = fresh_wire_2187[ 12 ];
	assign fresh_wire_2190[ 13 ] = fresh_wire_2187[ 13 ];
	assign fresh_wire_2190[ 14 ] = fresh_wire_2187[ 14 ];
	assign fresh_wire_2190[ 15 ] = fresh_wire_2187[ 15 ];
	assign fresh_wire_2190[ 16 ] = fresh_wire_2187[ 16 ];
	assign fresh_wire_2191[ 0 ] = fresh_wire_2189[ 0 ];
	assign fresh_wire_2191[ 1 ] = fresh_wire_2189[ 1 ];
	assign fresh_wire_2191[ 2 ] = fresh_wire_2189[ 2 ];
	assign fresh_wire_2191[ 3 ] = fresh_wire_2189[ 3 ];
	assign fresh_wire_2191[ 4 ] = fresh_wire_2189[ 4 ];
	assign fresh_wire_2191[ 5 ] = fresh_wire_2189[ 5 ];
	assign fresh_wire_2191[ 6 ] = fresh_wire_2189[ 6 ];
	assign fresh_wire_2191[ 7 ] = fresh_wire_2189[ 7 ];
	assign fresh_wire_2191[ 8 ] = fresh_wire_2189[ 8 ];
	assign fresh_wire_2191[ 9 ] = fresh_wire_2189[ 9 ];
	assign fresh_wire_2191[ 10 ] = fresh_wire_2189[ 10 ];
	assign fresh_wire_2191[ 11 ] = fresh_wire_2189[ 11 ];
	assign fresh_wire_2191[ 12 ] = fresh_wire_2189[ 12 ];
	assign fresh_wire_2191[ 13 ] = fresh_wire_2189[ 13 ];
	assign fresh_wire_2191[ 14 ] = fresh_wire_2189[ 14 ];
	assign fresh_wire_2191[ 15 ] = fresh_wire_2189[ 15 ];
	assign fresh_wire_2191[ 16 ] = fresh_wire_2189[ 16 ];
	assign fresh_wire_2193[ 0 ] = fresh_wire_2192[ 0 ];
	assign fresh_wire_2193[ 1 ] = fresh_wire_2192[ 1 ];
	assign fresh_wire_2193[ 2 ] = fresh_wire_2192[ 2 ];
	assign fresh_wire_2193[ 3 ] = fresh_wire_2192[ 3 ];
	assign fresh_wire_2193[ 4 ] = fresh_wire_2192[ 4 ];
	assign fresh_wire_2193[ 5 ] = fresh_wire_2192[ 5 ];
	assign fresh_wire_2193[ 6 ] = fresh_wire_2192[ 6 ];
	assign fresh_wire_2193[ 7 ] = fresh_wire_2192[ 7 ];
	assign fresh_wire_2193[ 8 ] = fresh_wire_2192[ 8 ];
	assign fresh_wire_2193[ 9 ] = fresh_wire_2192[ 9 ];
	assign fresh_wire_2193[ 10 ] = fresh_wire_2192[ 10 ];
	assign fresh_wire_2193[ 11 ] = fresh_wire_2192[ 11 ];
	assign fresh_wire_2193[ 12 ] = fresh_wire_2192[ 12 ];
	assign fresh_wire_2193[ 13 ] = fresh_wire_2192[ 13 ];
	assign fresh_wire_2193[ 14 ] = fresh_wire_2192[ 14 ];
	assign fresh_wire_2193[ 15 ] = fresh_wire_2192[ 15 ];
	assign fresh_wire_2193[ 16 ] = fresh_wire_2192[ 16 ];
	assign fresh_wire_2194[ 0 ] = fresh_wire_2296[ 0 ];
	assign fresh_wire_2194[ 1 ] = fresh_wire_2296[ 1 ];
	assign fresh_wire_2194[ 2 ] = fresh_wire_2296[ 2 ];
	assign fresh_wire_2194[ 3 ] = fresh_wire_2296[ 3 ];
	assign fresh_wire_2194[ 4 ] = fresh_wire_2296[ 4 ];
	assign fresh_wire_2194[ 5 ] = fresh_wire_2296[ 5 ];
	assign fresh_wire_2194[ 6 ] = fresh_wire_2296[ 6 ];
	assign fresh_wire_2194[ 7 ] = fresh_wire_2296[ 7 ];
	assign fresh_wire_2194[ 8 ] = fresh_wire_2296[ 8 ];
	assign fresh_wire_2194[ 9 ] = fresh_wire_2296[ 9 ];
	assign fresh_wire_2194[ 10 ] = fresh_wire_2296[ 10 ];
	assign fresh_wire_2194[ 11 ] = fresh_wire_2296[ 11 ];
	assign fresh_wire_2194[ 12 ] = fresh_wire_2296[ 12 ];
	assign fresh_wire_2194[ 13 ] = fresh_wire_2296[ 13 ];
	assign fresh_wire_2194[ 14 ] = fresh_wire_2296[ 14 ];
	assign fresh_wire_2194[ 15 ] = fresh_wire_2296[ 15 ];
	assign fresh_wire_2194[ 16 ] = fresh_wire_2296[ 16 ];
	assign fresh_wire_2196[ 0 ] = fresh_wire_2195[ 0 ];
	assign fresh_wire_2196[ 1 ] = fresh_wire_2195[ 1 ];
	assign fresh_wire_2196[ 2 ] = fresh_wire_2195[ 2 ];
	assign fresh_wire_2196[ 3 ] = fresh_wire_2195[ 3 ];
	assign fresh_wire_2196[ 4 ] = fresh_wire_2195[ 4 ];
	assign fresh_wire_2196[ 5 ] = fresh_wire_2195[ 5 ];
	assign fresh_wire_2196[ 6 ] = fresh_wire_2195[ 6 ];
	assign fresh_wire_2196[ 7 ] = fresh_wire_2195[ 7 ];
	assign fresh_wire_2196[ 8 ] = fresh_wire_2195[ 8 ];
	assign fresh_wire_2196[ 9 ] = fresh_wire_2195[ 9 ];
	assign fresh_wire_2196[ 10 ] = fresh_wire_2195[ 10 ];
	assign fresh_wire_2196[ 11 ] = fresh_wire_2195[ 11 ];
	assign fresh_wire_2196[ 12 ] = fresh_wire_2195[ 12 ];
	assign fresh_wire_2196[ 13 ] = fresh_wire_2195[ 13 ];
	assign fresh_wire_2196[ 14 ] = fresh_wire_2195[ 14 ];
	assign fresh_wire_2196[ 15 ] = fresh_wire_2195[ 15 ];
	assign fresh_wire_2198[ 0 ] = fresh_wire_2111[ 0 ];
	assign fresh_wire_2198[ 1 ] = fresh_wire_2111[ 1 ];
	assign fresh_wire_2198[ 2 ] = fresh_wire_2111[ 2 ];
	assign fresh_wire_2198[ 3 ] = fresh_wire_2111[ 3 ];
	assign fresh_wire_2198[ 4 ] = fresh_wire_2111[ 4 ];
	assign fresh_wire_2198[ 5 ] = fresh_wire_2111[ 5 ];
	assign fresh_wire_2198[ 6 ] = fresh_wire_2111[ 6 ];
	assign fresh_wire_2198[ 7 ] = fresh_wire_2111[ 7 ];
	assign fresh_wire_2198[ 8 ] = fresh_wire_2111[ 8 ];
	assign fresh_wire_2198[ 9 ] = fresh_wire_2111[ 9 ];
	assign fresh_wire_2198[ 10 ] = fresh_wire_2111[ 10 ];
	assign fresh_wire_2198[ 11 ] = fresh_wire_2111[ 11 ];
	assign fresh_wire_2198[ 12 ] = fresh_wire_2111[ 12 ];
	assign fresh_wire_2198[ 13 ] = fresh_wire_2111[ 13 ];
	assign fresh_wire_2198[ 14 ] = fresh_wire_2111[ 14 ];
	assign fresh_wire_2198[ 15 ] = fresh_wire_2111[ 15 ];
	assign fresh_wire_2200[ 0 ] = fresh_wire_2197[ 0 ];
	assign fresh_wire_2200[ 1 ] = fresh_wire_2197[ 1 ];
	assign fresh_wire_2200[ 2 ] = fresh_wire_2197[ 2 ];
	assign fresh_wire_2200[ 3 ] = fresh_wire_2197[ 3 ];
	assign fresh_wire_2200[ 4 ] = fresh_wire_2197[ 4 ];
	assign fresh_wire_2200[ 5 ] = fresh_wire_2197[ 5 ];
	assign fresh_wire_2200[ 6 ] = fresh_wire_2197[ 6 ];
	assign fresh_wire_2200[ 7 ] = fresh_wire_2197[ 7 ];
	assign fresh_wire_2200[ 8 ] = fresh_wire_2197[ 8 ];
	assign fresh_wire_2200[ 9 ] = fresh_wire_2197[ 9 ];
	assign fresh_wire_2200[ 10 ] = fresh_wire_2197[ 10 ];
	assign fresh_wire_2200[ 11 ] = fresh_wire_2197[ 11 ];
	assign fresh_wire_2200[ 12 ] = fresh_wire_2197[ 12 ];
	assign fresh_wire_2200[ 13 ] = fresh_wire_2197[ 13 ];
	assign fresh_wire_2200[ 14 ] = fresh_wire_2197[ 14 ];
	assign fresh_wire_2200[ 15 ] = fresh_wire_2197[ 15 ];
	assign fresh_wire_2200[ 16 ] = fresh_wire_2197[ 16 ];
	assign fresh_wire_2201[ 0 ] = fresh_wire_2199[ 0 ];
	assign fresh_wire_2201[ 1 ] = fresh_wire_2199[ 1 ];
	assign fresh_wire_2201[ 2 ] = fresh_wire_2199[ 2 ];
	assign fresh_wire_2201[ 3 ] = fresh_wire_2199[ 3 ];
	assign fresh_wire_2201[ 4 ] = fresh_wire_2199[ 4 ];
	assign fresh_wire_2201[ 5 ] = fresh_wire_2199[ 5 ];
	assign fresh_wire_2201[ 6 ] = fresh_wire_2199[ 6 ];
	assign fresh_wire_2201[ 7 ] = fresh_wire_2199[ 7 ];
	assign fresh_wire_2201[ 8 ] = fresh_wire_2199[ 8 ];
	assign fresh_wire_2201[ 9 ] = fresh_wire_2199[ 9 ];
	assign fresh_wire_2201[ 10 ] = fresh_wire_2199[ 10 ];
	assign fresh_wire_2201[ 11 ] = fresh_wire_2199[ 11 ];
	assign fresh_wire_2201[ 12 ] = fresh_wire_2199[ 12 ];
	assign fresh_wire_2201[ 13 ] = fresh_wire_2199[ 13 ];
	assign fresh_wire_2201[ 14 ] = fresh_wire_2199[ 14 ];
	assign fresh_wire_2201[ 15 ] = fresh_wire_2199[ 15 ];
	assign fresh_wire_2201[ 16 ] = fresh_wire_2199[ 16 ];
	assign fresh_wire_2203[ 0 ] = fresh_wire_2202[ 0 ];
	assign fresh_wire_2203[ 1 ] = fresh_wire_2202[ 1 ];
	assign fresh_wire_2203[ 2 ] = fresh_wire_2202[ 2 ];
	assign fresh_wire_2203[ 3 ] = fresh_wire_2202[ 3 ];
	assign fresh_wire_2203[ 4 ] = fresh_wire_2202[ 4 ];
	assign fresh_wire_2203[ 5 ] = fresh_wire_2202[ 5 ];
	assign fresh_wire_2203[ 6 ] = fresh_wire_2202[ 6 ];
	assign fresh_wire_2203[ 7 ] = fresh_wire_2202[ 7 ];
	assign fresh_wire_2203[ 8 ] = fresh_wire_2202[ 8 ];
	assign fresh_wire_2203[ 9 ] = fresh_wire_2202[ 9 ];
	assign fresh_wire_2203[ 10 ] = fresh_wire_2202[ 10 ];
	assign fresh_wire_2203[ 11 ] = fresh_wire_2202[ 11 ];
	assign fresh_wire_2203[ 12 ] = fresh_wire_2202[ 12 ];
	assign fresh_wire_2203[ 13 ] = fresh_wire_2202[ 13 ];
	assign fresh_wire_2203[ 14 ] = fresh_wire_2202[ 14 ];
	assign fresh_wire_2203[ 15 ] = fresh_wire_2202[ 15 ];
	assign fresh_wire_2203[ 16 ] = fresh_wire_2202[ 16 ];
	assign fresh_wire_2204[ 0 ] = fresh_wire_2297[ 0 ];
	assign fresh_wire_2204[ 1 ] = fresh_wire_2297[ 1 ];
	assign fresh_wire_2204[ 2 ] = fresh_wire_2297[ 2 ];
	assign fresh_wire_2204[ 3 ] = fresh_wire_2297[ 3 ];
	assign fresh_wire_2204[ 4 ] = fresh_wire_2297[ 4 ];
	assign fresh_wire_2204[ 5 ] = fresh_wire_2297[ 5 ];
	assign fresh_wire_2204[ 6 ] = fresh_wire_2297[ 6 ];
	assign fresh_wire_2204[ 7 ] = fresh_wire_2297[ 7 ];
	assign fresh_wire_2204[ 8 ] = fresh_wire_2297[ 8 ];
	assign fresh_wire_2204[ 9 ] = fresh_wire_2297[ 9 ];
	assign fresh_wire_2204[ 10 ] = fresh_wire_2297[ 10 ];
	assign fresh_wire_2204[ 11 ] = fresh_wire_2297[ 11 ];
	assign fresh_wire_2204[ 12 ] = fresh_wire_2297[ 12 ];
	assign fresh_wire_2204[ 13 ] = fresh_wire_2297[ 13 ];
	assign fresh_wire_2204[ 14 ] = fresh_wire_2297[ 14 ];
	assign fresh_wire_2204[ 15 ] = fresh_wire_2297[ 15 ];
	assign fresh_wire_2204[ 16 ] = fresh_wire_2297[ 16 ];
	assign fresh_wire_2206[ 0 ] = fresh_wire_2205[ 0 ];
	assign fresh_wire_2206[ 1 ] = fresh_wire_2205[ 1 ];
	assign fresh_wire_2206[ 2 ] = fresh_wire_2205[ 2 ];
	assign fresh_wire_2206[ 3 ] = fresh_wire_2205[ 3 ];
	assign fresh_wire_2206[ 4 ] = fresh_wire_2205[ 4 ];
	assign fresh_wire_2206[ 5 ] = fresh_wire_2205[ 5 ];
	assign fresh_wire_2206[ 6 ] = fresh_wire_2205[ 6 ];
	assign fresh_wire_2206[ 7 ] = fresh_wire_2205[ 7 ];
	assign fresh_wire_2206[ 8 ] = fresh_wire_2205[ 8 ];
	assign fresh_wire_2206[ 9 ] = fresh_wire_2205[ 9 ];
	assign fresh_wire_2206[ 10 ] = fresh_wire_2205[ 10 ];
	assign fresh_wire_2206[ 11 ] = fresh_wire_2205[ 11 ];
	assign fresh_wire_2206[ 12 ] = fresh_wire_2205[ 12 ];
	assign fresh_wire_2206[ 13 ] = fresh_wire_2205[ 13 ];
	assign fresh_wire_2206[ 14 ] = fresh_wire_2205[ 14 ];
	assign fresh_wire_2206[ 15 ] = fresh_wire_2205[ 15 ];
	assign fresh_wire_2208[ 0 ] = fresh_wire_2106[ 0 ];
	assign fresh_wire_2208[ 1 ] = fresh_wire_2106[ 1 ];
	assign fresh_wire_2208[ 2 ] = fresh_wire_2106[ 2 ];
	assign fresh_wire_2208[ 3 ] = fresh_wire_2106[ 3 ];
	assign fresh_wire_2208[ 4 ] = fresh_wire_2106[ 4 ];
	assign fresh_wire_2208[ 5 ] = fresh_wire_2106[ 5 ];
	assign fresh_wire_2208[ 6 ] = fresh_wire_2106[ 6 ];
	assign fresh_wire_2208[ 7 ] = fresh_wire_2106[ 7 ];
	assign fresh_wire_2208[ 8 ] = fresh_wire_2106[ 8 ];
	assign fresh_wire_2208[ 9 ] = fresh_wire_2106[ 9 ];
	assign fresh_wire_2208[ 10 ] = fresh_wire_2106[ 10 ];
	assign fresh_wire_2208[ 11 ] = fresh_wire_2106[ 11 ];
	assign fresh_wire_2208[ 12 ] = fresh_wire_2106[ 12 ];
	assign fresh_wire_2208[ 13 ] = fresh_wire_2106[ 13 ];
	assign fresh_wire_2208[ 14 ] = fresh_wire_2106[ 14 ];
	assign fresh_wire_2208[ 15 ] = fresh_wire_2106[ 15 ];
	assign fresh_wire_2210[ 0 ] = fresh_wire_2207[ 0 ];
	assign fresh_wire_2210[ 1 ] = fresh_wire_2207[ 1 ];
	assign fresh_wire_2210[ 2 ] = fresh_wire_2207[ 2 ];
	assign fresh_wire_2210[ 3 ] = fresh_wire_2207[ 3 ];
	assign fresh_wire_2210[ 4 ] = fresh_wire_2207[ 4 ];
	assign fresh_wire_2210[ 5 ] = fresh_wire_2207[ 5 ];
	assign fresh_wire_2210[ 6 ] = fresh_wire_2207[ 6 ];
	assign fresh_wire_2210[ 7 ] = fresh_wire_2207[ 7 ];
	assign fresh_wire_2210[ 8 ] = fresh_wire_2207[ 8 ];
	assign fresh_wire_2210[ 9 ] = fresh_wire_2207[ 9 ];
	assign fresh_wire_2210[ 10 ] = fresh_wire_2207[ 10 ];
	assign fresh_wire_2210[ 11 ] = fresh_wire_2207[ 11 ];
	assign fresh_wire_2210[ 12 ] = fresh_wire_2207[ 12 ];
	assign fresh_wire_2210[ 13 ] = fresh_wire_2207[ 13 ];
	assign fresh_wire_2210[ 14 ] = fresh_wire_2207[ 14 ];
	assign fresh_wire_2210[ 15 ] = fresh_wire_2207[ 15 ];
	assign fresh_wire_2210[ 16 ] = fresh_wire_2207[ 16 ];
	assign fresh_wire_2211[ 0 ] = fresh_wire_2209[ 0 ];
	assign fresh_wire_2211[ 1 ] = fresh_wire_2209[ 1 ];
	assign fresh_wire_2211[ 2 ] = fresh_wire_2209[ 2 ];
	assign fresh_wire_2211[ 3 ] = fresh_wire_2209[ 3 ];
	assign fresh_wire_2211[ 4 ] = fresh_wire_2209[ 4 ];
	assign fresh_wire_2211[ 5 ] = fresh_wire_2209[ 5 ];
	assign fresh_wire_2211[ 6 ] = fresh_wire_2209[ 6 ];
	assign fresh_wire_2211[ 7 ] = fresh_wire_2209[ 7 ];
	assign fresh_wire_2211[ 8 ] = fresh_wire_2209[ 8 ];
	assign fresh_wire_2211[ 9 ] = fresh_wire_2209[ 9 ];
	assign fresh_wire_2211[ 10 ] = fresh_wire_2209[ 10 ];
	assign fresh_wire_2211[ 11 ] = fresh_wire_2209[ 11 ];
	assign fresh_wire_2211[ 12 ] = fresh_wire_2209[ 12 ];
	assign fresh_wire_2211[ 13 ] = fresh_wire_2209[ 13 ];
	assign fresh_wire_2211[ 14 ] = fresh_wire_2209[ 14 ];
	assign fresh_wire_2211[ 15 ] = fresh_wire_2209[ 15 ];
	assign fresh_wire_2211[ 16 ] = fresh_wire_2209[ 16 ];
	assign fresh_wire_2213[ 0 ] = fresh_wire_2212[ 0 ];
	assign fresh_wire_2213[ 1 ] = fresh_wire_2212[ 1 ];
	assign fresh_wire_2213[ 2 ] = fresh_wire_2212[ 2 ];
	assign fresh_wire_2213[ 3 ] = fresh_wire_2212[ 3 ];
	assign fresh_wire_2213[ 4 ] = fresh_wire_2212[ 4 ];
	assign fresh_wire_2213[ 5 ] = fresh_wire_2212[ 5 ];
	assign fresh_wire_2213[ 6 ] = fresh_wire_2212[ 6 ];
	assign fresh_wire_2213[ 7 ] = fresh_wire_2212[ 7 ];
	assign fresh_wire_2213[ 8 ] = fresh_wire_2212[ 8 ];
	assign fresh_wire_2213[ 9 ] = fresh_wire_2212[ 9 ];
	assign fresh_wire_2213[ 10 ] = fresh_wire_2212[ 10 ];
	assign fresh_wire_2213[ 11 ] = fresh_wire_2212[ 11 ];
	assign fresh_wire_2213[ 12 ] = fresh_wire_2212[ 12 ];
	assign fresh_wire_2213[ 13 ] = fresh_wire_2212[ 13 ];
	assign fresh_wire_2213[ 14 ] = fresh_wire_2212[ 14 ];
	assign fresh_wire_2213[ 15 ] = fresh_wire_2212[ 15 ];
	assign fresh_wire_2213[ 16 ] = fresh_wire_2212[ 16 ];
	assign fresh_wire_2214[ 0 ] = fresh_wire_2298[ 0 ];
	assign fresh_wire_2214[ 1 ] = fresh_wire_2298[ 1 ];
	assign fresh_wire_2214[ 2 ] = fresh_wire_2298[ 2 ];
	assign fresh_wire_2214[ 3 ] = fresh_wire_2298[ 3 ];
	assign fresh_wire_2214[ 4 ] = fresh_wire_2298[ 4 ];
	assign fresh_wire_2214[ 5 ] = fresh_wire_2298[ 5 ];
	assign fresh_wire_2214[ 6 ] = fresh_wire_2298[ 6 ];
	assign fresh_wire_2214[ 7 ] = fresh_wire_2298[ 7 ];
	assign fresh_wire_2214[ 8 ] = fresh_wire_2298[ 8 ];
	assign fresh_wire_2214[ 9 ] = fresh_wire_2298[ 9 ];
	assign fresh_wire_2214[ 10 ] = fresh_wire_2298[ 10 ];
	assign fresh_wire_2214[ 11 ] = fresh_wire_2298[ 11 ];
	assign fresh_wire_2214[ 12 ] = fresh_wire_2298[ 12 ];
	assign fresh_wire_2214[ 13 ] = fresh_wire_2298[ 13 ];
	assign fresh_wire_2214[ 14 ] = fresh_wire_2298[ 14 ];
	assign fresh_wire_2214[ 15 ] = fresh_wire_2298[ 15 ];
	assign fresh_wire_2214[ 16 ] = fresh_wire_2298[ 16 ];
	assign fresh_wire_2216[ 0 ] = fresh_wire_2097[ 0 ];
	assign fresh_wire_2216[ 1 ] = fresh_wire_2097[ 1 ];
	assign fresh_wire_2216[ 2 ] = fresh_wire_2097[ 2 ];
	assign fresh_wire_2216[ 3 ] = fresh_wire_2097[ 3 ];
	assign fresh_wire_2216[ 4 ] = fresh_wire_2097[ 4 ];
	assign fresh_wire_2216[ 5 ] = fresh_wire_2097[ 5 ];
	assign fresh_wire_2216[ 6 ] = fresh_wire_2097[ 6 ];
	assign fresh_wire_2216[ 7 ] = fresh_wire_2097[ 7 ];
	assign fresh_wire_2216[ 8 ] = fresh_wire_2097[ 8 ];
	assign fresh_wire_2216[ 9 ] = fresh_wire_2097[ 9 ];
	assign fresh_wire_2216[ 10 ] = fresh_wire_2097[ 10 ];
	assign fresh_wire_2216[ 11 ] = fresh_wire_2097[ 11 ];
	assign fresh_wire_2216[ 12 ] = fresh_wire_2097[ 12 ];
	assign fresh_wire_2216[ 13 ] = fresh_wire_2097[ 13 ];
	assign fresh_wire_2216[ 14 ] = fresh_wire_2097[ 14 ];
	assign fresh_wire_2216[ 15 ] = fresh_wire_2097[ 15 ];
	assign fresh_wire_2216[ 16 ] = fresh_wire_2299[ 0 ];
	assign fresh_wire_2218[ 0 ] = fresh_wire_2217[ 0 ];
	assign fresh_wire_2218[ 1 ] = fresh_wire_2217[ 1 ];
	assign fresh_wire_2218[ 2 ] = fresh_wire_2217[ 2 ];
	assign fresh_wire_2218[ 3 ] = fresh_wire_2217[ 3 ];
	assign fresh_wire_2218[ 4 ] = fresh_wire_2217[ 4 ];
	assign fresh_wire_2218[ 5 ] = fresh_wire_2217[ 5 ];
	assign fresh_wire_2218[ 6 ] = fresh_wire_2217[ 6 ];
	assign fresh_wire_2218[ 7 ] = fresh_wire_2217[ 7 ];
	assign fresh_wire_2218[ 8 ] = fresh_wire_2217[ 8 ];
	assign fresh_wire_2218[ 9 ] = fresh_wire_2217[ 9 ];
	assign fresh_wire_2218[ 10 ] = fresh_wire_2217[ 10 ];
	assign fresh_wire_2218[ 11 ] = fresh_wire_2217[ 11 ];
	assign fresh_wire_2218[ 12 ] = fresh_wire_2217[ 12 ];
	assign fresh_wire_2218[ 13 ] = fresh_wire_2217[ 13 ];
	assign fresh_wire_2218[ 14 ] = fresh_wire_2217[ 14 ];
	assign fresh_wire_2218[ 15 ] = fresh_wire_2217[ 15 ];
	assign fresh_wire_2218[ 16 ] = fresh_wire_2217[ 16 ];
	assign fresh_wire_2218[ 17 ] = fresh_wire_2217[ 17 ];
	assign fresh_wire_2218[ 18 ] = fresh_wire_2217[ 18 ];
	assign fresh_wire_2218[ 19 ] = fresh_wire_2217[ 19 ];
	assign fresh_wire_2218[ 20 ] = fresh_wire_2217[ 20 ];
	assign fresh_wire_2218[ 21 ] = fresh_wire_2217[ 21 ];
	assign fresh_wire_2218[ 22 ] = fresh_wire_2217[ 22 ];
	assign fresh_wire_2218[ 23 ] = fresh_wire_2217[ 23 ];
	assign fresh_wire_2218[ 24 ] = fresh_wire_2217[ 24 ];
	assign fresh_wire_2218[ 25 ] = fresh_wire_2217[ 25 ];
	assign fresh_wire_2218[ 26 ] = fresh_wire_2217[ 26 ];
	assign fresh_wire_2218[ 27 ] = fresh_wire_2217[ 27 ];
	assign fresh_wire_2218[ 28 ] = fresh_wire_2217[ 28 ];
	assign fresh_wire_2218[ 29 ] = fresh_wire_2217[ 29 ];
	assign fresh_wire_2218[ 30 ] = fresh_wire_2217[ 30 ];
	assign fresh_wire_2218[ 31 ] = fresh_wire_2217[ 31 ];
	assign fresh_wire_2218[ 32 ] = fresh_wire_2217[ 32 ];
	assign fresh_wire_2218[ 33 ] = fresh_wire_2217[ 33 ];
	assign fresh_wire_2219[ 0 ] = fresh_wire_2300[ 0 ];
	assign fresh_wire_2219[ 1 ] = fresh_wire_2300[ 1 ];
	assign fresh_wire_2219[ 2 ] = fresh_wire_2300[ 2 ];
	assign fresh_wire_2219[ 3 ] = fresh_wire_2300[ 3 ];
	assign fresh_wire_2219[ 4 ] = fresh_wire_2300[ 4 ];
	assign fresh_wire_2219[ 5 ] = fresh_wire_2300[ 5 ];
	assign fresh_wire_2219[ 6 ] = fresh_wire_2300[ 6 ];
	assign fresh_wire_2219[ 7 ] = fresh_wire_2300[ 7 ];
	assign fresh_wire_2219[ 8 ] = fresh_wire_2300[ 8 ];
	assign fresh_wire_2219[ 9 ] = fresh_wire_2300[ 9 ];
	assign fresh_wire_2219[ 10 ] = fresh_wire_2300[ 10 ];
	assign fresh_wire_2219[ 11 ] = fresh_wire_2300[ 11 ];
	assign fresh_wire_2219[ 12 ] = fresh_wire_2300[ 12 ];
	assign fresh_wire_2219[ 13 ] = fresh_wire_2300[ 13 ];
	assign fresh_wire_2219[ 14 ] = fresh_wire_2300[ 14 ];
	assign fresh_wire_2219[ 15 ] = fresh_wire_2300[ 15 ];
	assign fresh_wire_2219[ 16 ] = fresh_wire_2300[ 16 ];
	assign fresh_wire_2219[ 17 ] = fresh_wire_2300[ 17 ];
	assign fresh_wire_2219[ 18 ] = fresh_wire_2300[ 18 ];
	assign fresh_wire_2219[ 19 ] = fresh_wire_2300[ 19 ];
	assign fresh_wire_2219[ 20 ] = fresh_wire_2300[ 20 ];
	assign fresh_wire_2219[ 21 ] = fresh_wire_2300[ 21 ];
	assign fresh_wire_2219[ 22 ] = fresh_wire_2300[ 22 ];
	assign fresh_wire_2219[ 23 ] = fresh_wire_2300[ 23 ];
	assign fresh_wire_2219[ 24 ] = fresh_wire_2300[ 24 ];
	assign fresh_wire_2219[ 25 ] = fresh_wire_2300[ 25 ];
	assign fresh_wire_2219[ 26 ] = fresh_wire_2300[ 26 ];
	assign fresh_wire_2219[ 27 ] = fresh_wire_2300[ 27 ];
	assign fresh_wire_2219[ 28 ] = fresh_wire_2300[ 28 ];
	assign fresh_wire_2219[ 29 ] = fresh_wire_2300[ 29 ];
	assign fresh_wire_2219[ 30 ] = fresh_wire_2300[ 30 ];
	assign fresh_wire_2219[ 31 ] = fresh_wire_2300[ 31 ];
	assign fresh_wire_2219[ 32 ] = fresh_wire_2300[ 32 ];
	assign fresh_wire_2219[ 33 ] = fresh_wire_2300[ 33 ];
	assign fresh_wire_2221[ 0 ] = fresh_wire_2097[ 0 ];
	assign fresh_wire_2221[ 1 ] = fresh_wire_2097[ 1 ];
	assign fresh_wire_2221[ 2 ] = fresh_wire_2097[ 2 ];
	assign fresh_wire_2221[ 3 ] = fresh_wire_2097[ 3 ];
	assign fresh_wire_2221[ 4 ] = fresh_wire_2097[ 4 ];
	assign fresh_wire_2221[ 5 ] = fresh_wire_2097[ 5 ];
	assign fresh_wire_2221[ 6 ] = fresh_wire_2097[ 6 ];
	assign fresh_wire_2221[ 7 ] = fresh_wire_2097[ 7 ];
	assign fresh_wire_2221[ 8 ] = fresh_wire_2097[ 8 ];
	assign fresh_wire_2221[ 9 ] = fresh_wire_2097[ 9 ];
	assign fresh_wire_2221[ 10 ] = fresh_wire_2097[ 10 ];
	assign fresh_wire_2221[ 11 ] = fresh_wire_2097[ 11 ];
	assign fresh_wire_2221[ 12 ] = fresh_wire_2097[ 12 ];
	assign fresh_wire_2221[ 13 ] = fresh_wire_2097[ 13 ];
	assign fresh_wire_2221[ 14 ] = fresh_wire_2097[ 14 ];
	assign fresh_wire_2221[ 15 ] = fresh_wire_2097[ 15 ];
	assign fresh_wire_2223[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_2224[ 0 ] = fresh_wire_2301[ 0 ];
	assign fresh_wire_2225[ 0 ] = fresh_wire_2222[ 0 ];
	assign fresh_wire_2225[ 1 ] = fresh_wire_2222[ 1 ];
	assign fresh_wire_2225[ 2 ] = fresh_wire_2222[ 2 ];
	assign fresh_wire_2225[ 3 ] = fresh_wire_2222[ 3 ];
	assign fresh_wire_2225[ 4 ] = fresh_wire_2222[ 4 ];
	assign fresh_wire_2225[ 5 ] = fresh_wire_2222[ 5 ];
	assign fresh_wire_2225[ 6 ] = fresh_wire_2222[ 6 ];
	assign fresh_wire_2225[ 7 ] = fresh_wire_2222[ 7 ];
	assign fresh_wire_2225[ 8 ] = fresh_wire_2222[ 8 ];
	assign fresh_wire_2225[ 9 ] = fresh_wire_2222[ 9 ];
	assign fresh_wire_2225[ 10 ] = fresh_wire_2222[ 10 ];
	assign fresh_wire_2225[ 11 ] = fresh_wire_2222[ 11 ];
	assign fresh_wire_2225[ 12 ] = fresh_wire_2222[ 12 ];
	assign fresh_wire_2225[ 13 ] = fresh_wire_2222[ 13 ];
	assign fresh_wire_2225[ 14 ] = fresh_wire_2222[ 14 ];
	assign fresh_wire_2225[ 15 ] = fresh_wire_2222[ 15 ];
	assign fresh_wire_2225[ 16 ] = fresh_wire_2302[ 0 ];
	assign fresh_wire_2227[ 0 ] = fresh_wire_2226[ 0 ];
	assign fresh_wire_2227[ 1 ] = fresh_wire_2226[ 1 ];
	assign fresh_wire_2227[ 2 ] = fresh_wire_2226[ 2 ];
	assign fresh_wire_2227[ 3 ] = fresh_wire_2226[ 3 ];
	assign fresh_wire_2227[ 4 ] = fresh_wire_2226[ 4 ];
	assign fresh_wire_2227[ 5 ] = fresh_wire_2226[ 5 ];
	assign fresh_wire_2227[ 6 ] = fresh_wire_2226[ 6 ];
	assign fresh_wire_2227[ 7 ] = fresh_wire_2226[ 7 ];
	assign fresh_wire_2227[ 8 ] = fresh_wire_2226[ 8 ];
	assign fresh_wire_2227[ 9 ] = fresh_wire_2226[ 9 ];
	assign fresh_wire_2227[ 10 ] = fresh_wire_2226[ 10 ];
	assign fresh_wire_2227[ 11 ] = fresh_wire_2226[ 11 ];
	assign fresh_wire_2227[ 12 ] = fresh_wire_2226[ 12 ];
	assign fresh_wire_2227[ 13 ] = fresh_wire_2226[ 13 ];
	assign fresh_wire_2227[ 14 ] = fresh_wire_2226[ 14 ];
	assign fresh_wire_2227[ 15 ] = fresh_wire_2226[ 15 ];
	assign fresh_wire_2227[ 16 ] = fresh_wire_2226[ 16 ];
	assign fresh_wire_2227[ 17 ] = fresh_wire_2226[ 17 ];
	assign fresh_wire_2227[ 18 ] = fresh_wire_2226[ 18 ];
	assign fresh_wire_2227[ 19 ] = fresh_wire_2226[ 19 ];
	assign fresh_wire_2227[ 20 ] = fresh_wire_2226[ 20 ];
	assign fresh_wire_2227[ 21 ] = fresh_wire_2226[ 21 ];
	assign fresh_wire_2227[ 22 ] = fresh_wire_2226[ 22 ];
	assign fresh_wire_2227[ 23 ] = fresh_wire_2226[ 23 ];
	assign fresh_wire_2227[ 24 ] = fresh_wire_2226[ 24 ];
	assign fresh_wire_2227[ 25 ] = fresh_wire_2226[ 25 ];
	assign fresh_wire_2227[ 26 ] = fresh_wire_2226[ 26 ];
	assign fresh_wire_2227[ 27 ] = fresh_wire_2226[ 27 ];
	assign fresh_wire_2227[ 28 ] = fresh_wire_2226[ 28 ];
	assign fresh_wire_2227[ 29 ] = fresh_wire_2226[ 29 ];
	assign fresh_wire_2227[ 30 ] = fresh_wire_2226[ 30 ];
	assign fresh_wire_2227[ 31 ] = fresh_wire_2226[ 31 ];
	assign fresh_wire_2227[ 32 ] = fresh_wire_2226[ 32 ];
	assign fresh_wire_2227[ 33 ] = fresh_wire_2226[ 33 ];
	assign fresh_wire_2228[ 0 ] = fresh_wire_2303[ 0 ];
	assign fresh_wire_2228[ 1 ] = fresh_wire_2303[ 1 ];
	assign fresh_wire_2228[ 2 ] = fresh_wire_2303[ 2 ];
	assign fresh_wire_2228[ 3 ] = fresh_wire_2303[ 3 ];
	assign fresh_wire_2228[ 4 ] = fresh_wire_2303[ 4 ];
	assign fresh_wire_2228[ 5 ] = fresh_wire_2303[ 5 ];
	assign fresh_wire_2228[ 6 ] = fresh_wire_2303[ 6 ];
	assign fresh_wire_2228[ 7 ] = fresh_wire_2303[ 7 ];
	assign fresh_wire_2228[ 8 ] = fresh_wire_2303[ 8 ];
	assign fresh_wire_2228[ 9 ] = fresh_wire_2303[ 9 ];
	assign fresh_wire_2228[ 10 ] = fresh_wire_2303[ 10 ];
	assign fresh_wire_2228[ 11 ] = fresh_wire_2303[ 11 ];
	assign fresh_wire_2228[ 12 ] = fresh_wire_2303[ 12 ];
	assign fresh_wire_2228[ 13 ] = fresh_wire_2303[ 13 ];
	assign fresh_wire_2228[ 14 ] = fresh_wire_2303[ 14 ];
	assign fresh_wire_2228[ 15 ] = fresh_wire_2303[ 15 ];
	assign fresh_wire_2228[ 16 ] = fresh_wire_2303[ 16 ];
	assign fresh_wire_2228[ 17 ] = fresh_wire_2303[ 17 ];
	assign fresh_wire_2228[ 18 ] = fresh_wire_2303[ 18 ];
	assign fresh_wire_2228[ 19 ] = fresh_wire_2303[ 19 ];
	assign fresh_wire_2228[ 20 ] = fresh_wire_2303[ 20 ];
	assign fresh_wire_2228[ 21 ] = fresh_wire_2303[ 21 ];
	assign fresh_wire_2228[ 22 ] = fresh_wire_2303[ 22 ];
	assign fresh_wire_2228[ 23 ] = fresh_wire_2303[ 23 ];
	assign fresh_wire_2228[ 24 ] = fresh_wire_2303[ 24 ];
	assign fresh_wire_2228[ 25 ] = fresh_wire_2303[ 25 ];
	assign fresh_wire_2228[ 26 ] = fresh_wire_2303[ 26 ];
	assign fresh_wire_2228[ 27 ] = fresh_wire_2303[ 27 ];
	assign fresh_wire_2228[ 28 ] = fresh_wire_2303[ 28 ];
	assign fresh_wire_2228[ 29 ] = fresh_wire_2303[ 29 ];
	assign fresh_wire_2228[ 30 ] = fresh_wire_2303[ 30 ];
	assign fresh_wire_2228[ 31 ] = fresh_wire_2303[ 31 ];
	assign fresh_wire_2228[ 32 ] = fresh_wire_2303[ 32 ];
	assign fresh_wire_2228[ 33 ] = fresh_wire_2303[ 33 ];
	assign fresh_wire_2230[ 0 ] = fresh_wire_2100[ 0 ];
	assign fresh_wire_2230[ 1 ] = fresh_wire_2100[ 1 ];
	assign fresh_wire_2230[ 2 ] = fresh_wire_2100[ 2 ];
	assign fresh_wire_2230[ 3 ] = fresh_wire_2100[ 3 ];
	assign fresh_wire_2230[ 4 ] = fresh_wire_2100[ 4 ];
	assign fresh_wire_2230[ 5 ] = fresh_wire_2100[ 5 ];
	assign fresh_wire_2230[ 6 ] = fresh_wire_2100[ 6 ];
	assign fresh_wire_2230[ 7 ] = fresh_wire_2100[ 7 ];
	assign fresh_wire_2230[ 8 ] = fresh_wire_2100[ 8 ];
	assign fresh_wire_2230[ 9 ] = fresh_wire_2100[ 9 ];
	assign fresh_wire_2230[ 10 ] = fresh_wire_2100[ 10 ];
	assign fresh_wire_2230[ 11 ] = fresh_wire_2100[ 11 ];
	assign fresh_wire_2230[ 12 ] = fresh_wire_2100[ 12 ];
	assign fresh_wire_2230[ 13 ] = fresh_wire_2100[ 13 ];
	assign fresh_wire_2230[ 14 ] = fresh_wire_2100[ 14 ];
	assign fresh_wire_2230[ 15 ] = fresh_wire_2100[ 15 ];
	assign fresh_wire_2232[ 0 ] = fresh_wire_2[ 0 ];
	assign fresh_wire_2233[ 0 ] = fresh_wire_2304[ 0 ];
	assign fresh_wire_2234[ 0 ] = fresh_wire_2231[ 0 ];
	assign fresh_wire_2234[ 1 ] = fresh_wire_2231[ 1 ];
	assign fresh_wire_2234[ 2 ] = fresh_wire_2231[ 2 ];
	assign fresh_wire_2234[ 3 ] = fresh_wire_2231[ 3 ];
	assign fresh_wire_2234[ 4 ] = fresh_wire_2231[ 4 ];
	assign fresh_wire_2234[ 5 ] = fresh_wire_2231[ 5 ];
	assign fresh_wire_2234[ 6 ] = fresh_wire_2231[ 6 ];
	assign fresh_wire_2234[ 7 ] = fresh_wire_2231[ 7 ];
	assign fresh_wire_2234[ 8 ] = fresh_wire_2231[ 8 ];
	assign fresh_wire_2234[ 9 ] = fresh_wire_2231[ 9 ];
	assign fresh_wire_2234[ 10 ] = fresh_wire_2231[ 10 ];
	assign fresh_wire_2234[ 11 ] = fresh_wire_2231[ 11 ];
	assign fresh_wire_2234[ 12 ] = fresh_wire_2231[ 12 ];
	assign fresh_wire_2234[ 13 ] = fresh_wire_2231[ 13 ];
	assign fresh_wire_2234[ 14 ] = fresh_wire_2231[ 14 ];
	assign fresh_wire_2234[ 15 ] = fresh_wire_2231[ 15 ];
	assign fresh_wire_2234[ 16 ] = fresh_wire_2305[ 0 ];
	assign fresh_wire_2236[ 0 ] = fresh_wire_2235[ 0 ];
	assign fresh_wire_2236[ 1 ] = fresh_wire_2235[ 1 ];
	assign fresh_wire_2236[ 2 ] = fresh_wire_2235[ 2 ];
	assign fresh_wire_2236[ 3 ] = fresh_wire_2235[ 3 ];
	assign fresh_wire_2236[ 4 ] = fresh_wire_2235[ 4 ];
	assign fresh_wire_2236[ 5 ] = fresh_wire_2235[ 5 ];
	assign fresh_wire_2236[ 6 ] = fresh_wire_2235[ 6 ];
	assign fresh_wire_2236[ 7 ] = fresh_wire_2235[ 7 ];
	assign fresh_wire_2236[ 8 ] = fresh_wire_2235[ 8 ];
	assign fresh_wire_2236[ 9 ] = fresh_wire_2235[ 9 ];
	assign fresh_wire_2236[ 10 ] = fresh_wire_2235[ 10 ];
	assign fresh_wire_2236[ 11 ] = fresh_wire_2235[ 11 ];
	assign fresh_wire_2236[ 12 ] = fresh_wire_2235[ 12 ];
	assign fresh_wire_2236[ 13 ] = fresh_wire_2235[ 13 ];
	assign fresh_wire_2236[ 14 ] = fresh_wire_2235[ 14 ];
	assign fresh_wire_2236[ 15 ] = fresh_wire_2235[ 15 ];
	assign fresh_wire_2236[ 16 ] = fresh_wire_2235[ 16 ];
	assign fresh_wire_2236[ 17 ] = fresh_wire_2235[ 17 ];
	assign fresh_wire_2236[ 18 ] = fresh_wire_2235[ 18 ];
	assign fresh_wire_2236[ 19 ] = fresh_wire_2235[ 19 ];
	assign fresh_wire_2236[ 20 ] = fresh_wire_2235[ 20 ];
	assign fresh_wire_2236[ 21 ] = fresh_wire_2235[ 21 ];
	assign fresh_wire_2236[ 22 ] = fresh_wire_2235[ 22 ];
	assign fresh_wire_2236[ 23 ] = fresh_wire_2235[ 23 ];
	assign fresh_wire_2236[ 24 ] = fresh_wire_2235[ 24 ];
	assign fresh_wire_2236[ 25 ] = fresh_wire_2235[ 25 ];
	assign fresh_wire_2236[ 26 ] = fresh_wire_2235[ 26 ];
	assign fresh_wire_2236[ 27 ] = fresh_wire_2235[ 27 ];
	assign fresh_wire_2236[ 28 ] = fresh_wire_2235[ 28 ];
	assign fresh_wire_2236[ 29 ] = fresh_wire_2235[ 29 ];
	assign fresh_wire_2236[ 30 ] = fresh_wire_2235[ 30 ];
	assign fresh_wire_2236[ 31 ] = fresh_wire_2235[ 31 ];
	assign fresh_wire_2236[ 32 ] = fresh_wire_2235[ 32 ];
	assign fresh_wire_2236[ 33 ] = fresh_wire_2235[ 33 ];
	assign fresh_wire_2237[ 0 ] = fresh_wire_2306[ 0 ];
	assign fresh_wire_2237[ 1 ] = fresh_wire_2306[ 1 ];
	assign fresh_wire_2237[ 2 ] = fresh_wire_2306[ 2 ];
	assign fresh_wire_2237[ 3 ] = fresh_wire_2306[ 3 ];
	assign fresh_wire_2237[ 4 ] = fresh_wire_2306[ 4 ];
	assign fresh_wire_2237[ 5 ] = fresh_wire_2306[ 5 ];
	assign fresh_wire_2237[ 6 ] = fresh_wire_2306[ 6 ];
	assign fresh_wire_2237[ 7 ] = fresh_wire_2306[ 7 ];
	assign fresh_wire_2237[ 8 ] = fresh_wire_2306[ 8 ];
	assign fresh_wire_2237[ 9 ] = fresh_wire_2306[ 9 ];
	assign fresh_wire_2237[ 10 ] = fresh_wire_2306[ 10 ];
	assign fresh_wire_2237[ 11 ] = fresh_wire_2306[ 11 ];
	assign fresh_wire_2237[ 12 ] = fresh_wire_2306[ 12 ];
	assign fresh_wire_2237[ 13 ] = fresh_wire_2306[ 13 ];
	assign fresh_wire_2237[ 14 ] = fresh_wire_2306[ 14 ];
	assign fresh_wire_2237[ 15 ] = fresh_wire_2306[ 15 ];
	assign fresh_wire_2237[ 16 ] = fresh_wire_2306[ 16 ];
	assign fresh_wire_2237[ 17 ] = fresh_wire_2306[ 17 ];
	assign fresh_wire_2237[ 18 ] = fresh_wire_2306[ 18 ];
	assign fresh_wire_2237[ 19 ] = fresh_wire_2306[ 19 ];
	assign fresh_wire_2237[ 20 ] = fresh_wire_2306[ 20 ];
	assign fresh_wire_2237[ 21 ] = fresh_wire_2306[ 21 ];
	assign fresh_wire_2237[ 22 ] = fresh_wire_2306[ 22 ];
	assign fresh_wire_2237[ 23 ] = fresh_wire_2306[ 23 ];
	assign fresh_wire_2237[ 24 ] = fresh_wire_2306[ 24 ];
	assign fresh_wire_2237[ 25 ] = fresh_wire_2306[ 25 ];
	assign fresh_wire_2237[ 26 ] = fresh_wire_2306[ 26 ];
	assign fresh_wire_2237[ 27 ] = fresh_wire_2306[ 27 ];
	assign fresh_wire_2237[ 28 ] = fresh_wire_2306[ 28 ];
	assign fresh_wire_2237[ 29 ] = fresh_wire_2306[ 29 ];
	assign fresh_wire_2237[ 30 ] = fresh_wire_2306[ 30 ];
	assign fresh_wire_2237[ 31 ] = fresh_wire_2306[ 31 ];
	assign fresh_wire_2237[ 32 ] = fresh_wire_2306[ 32 ];
	assign fresh_wire_2237[ 33 ] = fresh_wire_2306[ 33 ];
	assign fresh_wire_2239[ 0 ] = fresh_wire_2220[ 0 ];
	assign fresh_wire_2239[ 1 ] = fresh_wire_2220[ 1 ];
	assign fresh_wire_2239[ 2 ] = fresh_wire_2220[ 2 ];
	assign fresh_wire_2239[ 3 ] = fresh_wire_2220[ 3 ];
	assign fresh_wire_2239[ 4 ] = fresh_wire_2220[ 4 ];
	assign fresh_wire_2239[ 5 ] = fresh_wire_2220[ 5 ];
	assign fresh_wire_2239[ 6 ] = fresh_wire_2220[ 6 ];
	assign fresh_wire_2239[ 7 ] = fresh_wire_2220[ 7 ];
	assign fresh_wire_2239[ 8 ] = fresh_wire_2220[ 8 ];
	assign fresh_wire_2239[ 9 ] = fresh_wire_2220[ 9 ];
	assign fresh_wire_2239[ 10 ] = fresh_wire_2220[ 10 ];
	assign fresh_wire_2239[ 11 ] = fresh_wire_2220[ 11 ];
	assign fresh_wire_2239[ 12 ] = fresh_wire_2220[ 12 ];
	assign fresh_wire_2239[ 13 ] = fresh_wire_2220[ 13 ];
	assign fresh_wire_2239[ 14 ] = fresh_wire_2220[ 14 ];
	assign fresh_wire_2239[ 15 ] = fresh_wire_2220[ 15 ];
	assign fresh_wire_2241[ 0 ] = fresh_wire_2185[ 0 ];
	assign fresh_wire_2241[ 1 ] = fresh_wire_2185[ 1 ];
	assign fresh_wire_2241[ 2 ] = fresh_wire_2185[ 2 ];
	assign fresh_wire_2241[ 3 ] = fresh_wire_2185[ 3 ];
	assign fresh_wire_2241[ 4 ] = fresh_wire_2185[ 4 ];
	assign fresh_wire_2241[ 5 ] = fresh_wire_2185[ 5 ];
	assign fresh_wire_2241[ 6 ] = fresh_wire_2185[ 6 ];
	assign fresh_wire_2241[ 7 ] = fresh_wire_2185[ 7 ];
	assign fresh_wire_2241[ 8 ] = fresh_wire_2185[ 8 ];
	assign fresh_wire_2241[ 9 ] = fresh_wire_2185[ 9 ];
	assign fresh_wire_2241[ 10 ] = fresh_wire_2185[ 10 ];
	assign fresh_wire_2241[ 11 ] = fresh_wire_2185[ 11 ];
	assign fresh_wire_2241[ 12 ] = fresh_wire_2185[ 12 ];
	assign fresh_wire_2241[ 13 ] = fresh_wire_2185[ 13 ];
	assign fresh_wire_2241[ 14 ] = fresh_wire_2185[ 14 ];
	assign fresh_wire_2241[ 15 ] = fresh_wire_2185[ 15 ];
	assign fresh_wire_2243[ 0 ] = fresh_wire_2240[ 0 ];
	assign fresh_wire_2243[ 1 ] = fresh_wire_2240[ 1 ];
	assign fresh_wire_2243[ 2 ] = fresh_wire_2240[ 2 ];
	assign fresh_wire_2243[ 3 ] = fresh_wire_2240[ 3 ];
	assign fresh_wire_2243[ 4 ] = fresh_wire_2240[ 4 ];
	assign fresh_wire_2243[ 5 ] = fresh_wire_2240[ 5 ];
	assign fresh_wire_2243[ 6 ] = fresh_wire_2240[ 6 ];
	assign fresh_wire_2243[ 7 ] = fresh_wire_2240[ 7 ];
	assign fresh_wire_2243[ 8 ] = fresh_wire_2240[ 8 ];
	assign fresh_wire_2243[ 9 ] = fresh_wire_2240[ 9 ];
	assign fresh_wire_2243[ 10 ] = fresh_wire_2240[ 10 ];
	assign fresh_wire_2243[ 11 ] = fresh_wire_2240[ 11 ];
	assign fresh_wire_2243[ 12 ] = fresh_wire_2240[ 12 ];
	assign fresh_wire_2243[ 13 ] = fresh_wire_2240[ 13 ];
	assign fresh_wire_2243[ 14 ] = fresh_wire_2240[ 14 ];
	assign fresh_wire_2243[ 15 ] = fresh_wire_2240[ 15 ];
	assign fresh_wire_2243[ 16 ] = fresh_wire_2240[ 16 ];
	assign fresh_wire_2244[ 0 ] = fresh_wire_2242[ 0 ];
	assign fresh_wire_2244[ 1 ] = fresh_wire_2242[ 1 ];
	assign fresh_wire_2244[ 2 ] = fresh_wire_2242[ 2 ];
	assign fresh_wire_2244[ 3 ] = fresh_wire_2242[ 3 ];
	assign fresh_wire_2244[ 4 ] = fresh_wire_2242[ 4 ];
	assign fresh_wire_2244[ 5 ] = fresh_wire_2242[ 5 ];
	assign fresh_wire_2244[ 6 ] = fresh_wire_2242[ 6 ];
	assign fresh_wire_2244[ 7 ] = fresh_wire_2242[ 7 ];
	assign fresh_wire_2244[ 8 ] = fresh_wire_2242[ 8 ];
	assign fresh_wire_2244[ 9 ] = fresh_wire_2242[ 9 ];
	assign fresh_wire_2244[ 10 ] = fresh_wire_2242[ 10 ];
	assign fresh_wire_2244[ 11 ] = fresh_wire_2242[ 11 ];
	assign fresh_wire_2244[ 12 ] = fresh_wire_2242[ 12 ];
	assign fresh_wire_2244[ 13 ] = fresh_wire_2242[ 13 ];
	assign fresh_wire_2244[ 14 ] = fresh_wire_2242[ 14 ];
	assign fresh_wire_2244[ 15 ] = fresh_wire_2242[ 15 ];
	assign fresh_wire_2244[ 16 ] = fresh_wire_2242[ 16 ];
	assign fresh_wire_2246[ 0 ] = fresh_wire_2245[ 0 ];
	assign fresh_wire_2246[ 1 ] = fresh_wire_2245[ 1 ];
	assign fresh_wire_2246[ 2 ] = fresh_wire_2245[ 2 ];
	assign fresh_wire_2246[ 3 ] = fresh_wire_2245[ 3 ];
	assign fresh_wire_2246[ 4 ] = fresh_wire_2245[ 4 ];
	assign fresh_wire_2246[ 5 ] = fresh_wire_2245[ 5 ];
	assign fresh_wire_2246[ 6 ] = fresh_wire_2245[ 6 ];
	assign fresh_wire_2246[ 7 ] = fresh_wire_2245[ 7 ];
	assign fresh_wire_2246[ 8 ] = fresh_wire_2245[ 8 ];
	assign fresh_wire_2246[ 9 ] = fresh_wire_2245[ 9 ];
	assign fresh_wire_2246[ 10 ] = fresh_wire_2245[ 10 ];
	assign fresh_wire_2246[ 11 ] = fresh_wire_2245[ 11 ];
	assign fresh_wire_2246[ 12 ] = fresh_wire_2245[ 12 ];
	assign fresh_wire_2246[ 13 ] = fresh_wire_2245[ 13 ];
	assign fresh_wire_2246[ 14 ] = fresh_wire_2245[ 14 ];
	assign fresh_wire_2246[ 15 ] = fresh_wire_2245[ 15 ];
	assign fresh_wire_2246[ 16 ] = fresh_wire_2245[ 16 ];
	assign fresh_wire_2247[ 0 ] = fresh_wire_2307[ 0 ];
	assign fresh_wire_2247[ 1 ] = fresh_wire_2307[ 1 ];
	assign fresh_wire_2247[ 2 ] = fresh_wire_2307[ 2 ];
	assign fresh_wire_2247[ 3 ] = fresh_wire_2307[ 3 ];
	assign fresh_wire_2247[ 4 ] = fresh_wire_2307[ 4 ];
	assign fresh_wire_2247[ 5 ] = fresh_wire_2307[ 5 ];
	assign fresh_wire_2247[ 6 ] = fresh_wire_2307[ 6 ];
	assign fresh_wire_2247[ 7 ] = fresh_wire_2307[ 7 ];
	assign fresh_wire_2247[ 8 ] = fresh_wire_2307[ 8 ];
	assign fresh_wire_2247[ 9 ] = fresh_wire_2307[ 9 ];
	assign fresh_wire_2247[ 10 ] = fresh_wire_2307[ 10 ];
	assign fresh_wire_2247[ 11 ] = fresh_wire_2307[ 11 ];
	assign fresh_wire_2247[ 12 ] = fresh_wire_2307[ 12 ];
	assign fresh_wire_2247[ 13 ] = fresh_wire_2307[ 13 ];
	assign fresh_wire_2247[ 14 ] = fresh_wire_2307[ 14 ];
	assign fresh_wire_2247[ 15 ] = fresh_wire_2307[ 15 ];
	assign fresh_wire_2247[ 16 ] = fresh_wire_2307[ 16 ];
endmodule

