module CELL_TYPE_CONST #(parameter PARAM_WIDTH=1, parameter PARAM_INIT_VALUE=0) (output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT); assign PORT_ID_OUT = PARAM_INIT_VALUE;
endmodule

module CELL_TYPE_MUL #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT); assign PORT_ID_OUT = PORT_ID_IN0 * PORT_ID_IN1;
 endmodule

module CELL_TYPE_NOT #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT); assign PORT_ID_OUT = ~PORT_ID_IN;
 endmodule

module CELL_TYPE_ADD #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT);
   assign PORT_ID_OUT = PORT_ID_IN0 + PORT_ID_IN1;
 endmodule

module CELL_TYPE_SUB #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT);   assign PORT_ID_OUT = PORT_ID_IN0 - PORT_ID_IN1; endmodule

module CELL_TYPE_AND #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT);
   assign PORT_ID_OUT = PORT_ID_IN0 & PORT_ID_IN1;
endmodule

module CELL_TYPE_OR #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT);
   assign PORT_ID_OUT = PORT_ID_IN0 | PORT_ID_IN1;
endmodule

module CELL_TYPE_EQ #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [0 : 0] PORT_ID_OUT);
   assign PORT_ID_OUT = PORT_ID_IN0 == PORT_ID_IN1;
endmodule

module CELL_TYPE_ULT #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [0 : 0] PORT_ID_OUT); assign PORT_ID_OUT = PORT_ID_IN0 < PORT_ID_IN1;
 endmodule

module CELL_TYPE_UGE #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [0 : 0] PORT_ID_OUT); assign PORT_ID_OUT = PORT_ID_IN0 >= PORT_ID_IN1;
endmodule

 // CELL_TYPE_UGE
module CELL_TYPE_REG #(parameter PARAM_CLK_POSEDGE=1, parameter PARAM_INIT_VALUE=0, parameter PARAM_WIDTH=1)(input PORT_ID_CLK, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT);
   reg [PARAM_WIDTH - 1 : 0] data;
   initial begin
      data = PARAM_INIT_VALUE;
   end
   wire true_clk;
   assign true_clk = PARAM_CLK_POSEDGE ? PORT_ID_CLK : ~PORT_ID_CLK;
   always @(posedge true_clk) begin
      data <= PORT_ID_IN;
   end
   assign PORT_ID_OUT = data;
endmodule

module CELL_TYPE_REG_ARST #(parameter PARAM_CLK_POSEDGE=1, parameter PARAM_ARST_POSEDGE=1, parameter PARAM_INIT_VALUE=0, parameter PARAM_WIDTH=1)(input PORT_ID_ARST, input PORT_ID_CLK, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT);
   reg [PARAM_WIDTH - 1 : 0] data;
   initial begin
      data = PARAM_INIT_VALUE;
   end
   wire true_clk;
   assign true_clk = PARAM_CLK_POSEDGE ? PORT_ID_CLK : ~PORT_ID_CLK;
   wire true_rst;
   assign true_rst = PARAM_ARST_POSEDGE ? PORT_ID_ARST : ~PORT_ID_ARST;
   always @(posedge true_clk or posedge true_rst) begin
      if (true_rst) begin
         data <= PARAM_INIT_VALUE;
      end else begin
         data <= PORT_ID_IN;
      end
   end
   assign PORT_ID_OUT = data;
endmodule

 // CELL_TYPE_REG_ARST
module CELL_TYPE_MEM #(parameter PARAM_HAS_INIT=0, parameter PARAM_MEM_DEPTH=0, parameter PARAM_MEM_WIDTH=0)(input PORT_ID_CLK, input PORT_ID_WEN, input [$clog2(PARAM_MEM_DEPTH) - 1 : 0] PORT_ID_RADDR, input [$clog2(PARAM_MEM_DEPTH) - 1 : 0] PORT_ID_WADDR, input [PARAM_MEM_WIDTH - 1 : 0] PORT_ID_WDATA, output [PARAM_MEM_WIDTH - 1 : 0] PORT_ID_RDATA);
   reg [PARAM_MEM_WIDTH -  1 : 0] data_array [0 : PARAM_MEM_DEPTH - 1];
   always @(posedge PORT_ID_CLK) begin
      if (PORT_ID_WEN) begin
         data_array[PORT_ID_WADDR] = PORT_ID_WDATA;
      end
   end
   assign PORT_ID_RDATA = data_array[PORT_ID_RADDR];
endmodule

module CELL_TYPE_MUX #(parameter PARAM_WIDTH=1) (input PORT_ID_SEL, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN0, input [PARAM_WIDTH - 1 : 0] PORT_ID_IN1, output [PARAM_WIDTH - 1 : 0] PORT_ID_OUT);
   assign PORT_ID_OUT = PORT_ID_SEL ? PORT_ID_IN1 : PORT_ID_IN0;
 endmodule

module CELL_TYPE_ORR #(parameter PARAM_WIDTH=1) (input [PARAM_WIDTH - 1 : 0] PORT_ID_IN, output [0 : 0] PORT_ID_OUT); assign PORT_ID_OUT = |PORT_ID_IN;
 endmodule

module CELL_TYPE_PORT #(parameter PARAM_PORT_TYPE=0, parameter PARAM_OUT_WIDTH=1) (input [PARAM_OUT_WIDTH - 1 : 0] PORT_ID_IN, output [PARAM_OUT_WIDTH - 1 : 0] PORT_ID_OUT); assign PORT_ID_OUT = PORT_ID_IN;
 endmodule

module CELL_TYPE_ZEXT #(parameter PARAM_IN_WIDTH=1, parameter PARAM_OUT_WIDTH=1) (input [PARAM_IN_WIDTH - 1 : 0] PORT_ID_IN, output [PARAM_OUT_WIDTH - 1 : 0] PORT_ID_OUT); assign PORT_ID_OUT = {{(PARAM_OUT_WIDTH - PARAM_IN_WIDTH){1'b0}}, PORT_ID_IN};
 endmodule


module flat_module(	output [0 : 0] aux_div_pad,
	input [0 : 0] clk_ext_in,
	input [0 : 0] clk_in,
	input [31 : 0] config_addr_in,
	input [31 : 0] config_data_in,
	input [0 : 0] ext_cki,
	input [0 : 0] ext_cki_jm,
	input [0 : 0] ext_ckib,
	input [0 : 0] ext_ckib_jm,
	input [0 : 0] ext_frefn,
	input [0 : 0] ext_frefn_jm,
	input [0 : 0] ext_frefp,
	input [0 : 0] ext_frefp_jm,
	output [0 : 0] ffeed_pad,
	output [0 : 0] fout_div_pad,
	output [0 : 0] fref_off_pad,
	output [0 : 0] frefn_out_jm,
	output [0 : 0] frefp_out_jm,
	output [12 : 0] lf_out,
	output [3 : 0] mdllout_pad,
	input [0 : 0] pad_S0_T0_in,
	output [0 : 0] pad_S0_T0_out,
	input [0 : 0] pad_S0_T10_in,
	output [0 : 0] pad_S0_T10_out,
	input [0 : 0] pad_S0_T11_in,
	output [0 : 0] pad_S0_T11_out,
	input [0 : 0] pad_S0_T12_in,
	output [0 : 0] pad_S0_T12_out,
	input [0 : 0] pad_S0_T13_in,
	output [0 : 0] pad_S0_T13_out,
	input [0 : 0] pad_S0_T14_in,
	output [0 : 0] pad_S0_T14_out,
	input [0 : 0] pad_S0_T15_in,
	output [0 : 0] pad_S0_T15_out,
	input [0 : 0] pad_S0_T1_in,
	output [0 : 0] pad_S0_T1_out,
	input [0 : 0] pad_S0_T2_in,
	output [0 : 0] pad_S0_T2_out,
	input [0 : 0] pad_S0_T3_in,
	output [0 : 0] pad_S0_T3_out,
	input [0 : 0] pad_S0_T4_in,
	output [0 : 0] pad_S0_T4_out,
	input [0 : 0] pad_S0_T5_in,
	output [0 : 0] pad_S0_T5_out,
	input [0 : 0] pad_S0_T6_in,
	output [0 : 0] pad_S0_T6_out,
	input [0 : 0] pad_S0_T7_in,
	output [0 : 0] pad_S0_T7_out,
	input [0 : 0] pad_S0_T8_in,
	output [0 : 0] pad_S0_T8_out,
	input [0 : 0] pad_S0_T9_in,
	output [0 : 0] pad_S0_T9_out,
	input [0 : 0] pad_S1_T0_in,
	output [0 : 0] pad_S1_T0_out,
	input [0 : 0] pad_S1_T10_in,
	output [0 : 0] pad_S1_T10_out,
	input [0 : 0] pad_S1_T11_in,
	output [0 : 0] pad_S1_T11_out,
	input [0 : 0] pad_S1_T12_in,
	output [0 : 0] pad_S1_T12_out,
	input [0 : 0] pad_S1_T13_in,
	output [0 : 0] pad_S1_T13_out,
	input [0 : 0] pad_S1_T14_in,
	output [0 : 0] pad_S1_T14_out,
	input [0 : 0] pad_S1_T15_in,
	output [0 : 0] pad_S1_T15_out,
	input [0 : 0] pad_S1_T1_in,
	output [0 : 0] pad_S1_T1_out,
	input [0 : 0] pad_S1_T2_in,
	output [0 : 0] pad_S1_T2_out,
	input [0 : 0] pad_S1_T3_in,
	output [0 : 0] pad_S1_T3_out,
	input [0 : 0] pad_S1_T4_in,
	output [0 : 0] pad_S1_T4_out,
	input [0 : 0] pad_S1_T5_in,
	output [0 : 0] pad_S1_T5_out,
	input [0 : 0] pad_S1_T6_in,
	output [0 : 0] pad_S1_T6_out,
	input [0 : 0] pad_S1_T7_in,
	output [0 : 0] pad_S1_T7_out,
	input [0 : 0] pad_S1_T8_in,
	output [0 : 0] pad_S1_T8_out,
	input [0 : 0] pad_S1_T9_in,
	output [0 : 0] pad_S1_T9_out,
	input [0 : 0] pad_S2_T0_in,
	output [0 : 0] pad_S2_T0_out,
	input [0 : 0] pad_S2_T10_in,
	output [0 : 0] pad_S2_T10_out,
	input [0 : 0] pad_S2_T11_in,
	output [0 : 0] pad_S2_T11_out,
	input [0 : 0] pad_S2_T12_in,
	output [0 : 0] pad_S2_T12_out,
	input [0 : 0] pad_S2_T13_in,
	output [0 : 0] pad_S2_T13_out,
	input [0 : 0] pad_S2_T14_in,
	output [0 : 0] pad_S2_T14_out,
	input [0 : 0] pad_S2_T15_in,
	output [0 : 0] pad_S2_T15_out,
	input [0 : 0] pad_S2_T1_in,
	output [0 : 0] pad_S2_T1_out,
	input [0 : 0] pad_S2_T2_in,
	output [0 : 0] pad_S2_T2_out,
	input [0 : 0] pad_S2_T3_in,
	output [0 : 0] pad_S2_T3_out,
	input [0 : 0] pad_S2_T4_in,
	output [0 : 0] pad_S2_T4_out,
	input [0 : 0] pad_S2_T5_in,
	output [0 : 0] pad_S2_T5_out,
	input [0 : 0] pad_S2_T6_in,
	output [0 : 0] pad_S2_T6_out,
	input [0 : 0] pad_S2_T7_in,
	output [0 : 0] pad_S2_T7_out,
	input [0 : 0] pad_S2_T8_in,
	output [0 : 0] pad_S2_T8_out,
	input [0 : 0] pad_S2_T9_in,
	output [0 : 0] pad_S2_T9_out,
	input [0 : 0] pad_S3_T0_in,
	output [0 : 0] pad_S3_T0_out,
	input [0 : 0] pad_S3_T10_in,
	output [0 : 0] pad_S3_T10_out,
	input [0 : 0] pad_S3_T11_in,
	output [0 : 0] pad_S3_T11_out,
	input [0 : 0] pad_S3_T12_in,
	output [0 : 0] pad_S3_T12_out,
	input [0 : 0] pad_S3_T13_in,
	output [0 : 0] pad_S3_T13_out,
	input [0 : 0] pad_S3_T14_in,
	output [0 : 0] pad_S3_T14_out,
	input [0 : 0] pad_S3_T15_in,
	output [0 : 0] pad_S3_T15_out,
	input [0 : 0] pad_S3_T1_in,
	output [0 : 0] pad_S3_T1_out,
	input [0 : 0] pad_S3_T2_in,
	output [0 : 0] pad_S3_T2_out,
	input [0 : 0] pad_S3_T3_in,
	output [0 : 0] pad_S3_T3_out,
	input [0 : 0] pad_S3_T4_in,
	output [0 : 0] pad_S3_T4_out,
	input [0 : 0] pad_S3_T5_in,
	output [0 : 0] pad_S3_T5_out,
	input [0 : 0] pad_S3_T6_in,
	output [0 : 0] pad_S3_T6_out,
	input [0 : 0] pad_S3_T7_in,
	output [0 : 0] pad_S3_T7_out,
	input [0 : 0] pad_S3_T8_in,
	output [0 : 0] pad_S3_T8_out,
	input [0 : 0] pad_S3_T9_in,
	output [0 : 0] pad_S3_T9_out,
	input [0 : 0] reset_in,
	input [0 : 0] tck,
	input [0 : 0] tdi,
	output [0 : 0] tdo,
	input [0 : 0] tms,
	input [0 : 0] trst_n);

	wire [0 : 0] fresh_wire_0;
	wire [0 : 0] fresh_wire_1;
	wire [0 : 0] fresh_wire_2;
	wire [31 : 0] fresh_wire_3;
	wire [31 : 0] fresh_wire_4;
	wire [0 : 0] fresh_wire_5;
	wire [0 : 0] fresh_wire_6;
	wire [0 : 0] fresh_wire_7;
	wire [0 : 0] fresh_wire_8;
	wire [0 : 0] fresh_wire_9;
	wire [0 : 0] fresh_wire_10;
	wire [0 : 0] fresh_wire_11;
	wire [0 : 0] fresh_wire_12;
	wire [0 : 0] fresh_wire_13;
	wire [0 : 0] fresh_wire_14;
	wire [0 : 0] fresh_wire_15;
	wire [0 : 0] fresh_wire_16;
	wire [0 : 0] fresh_wire_17;
	wire [12 : 0] fresh_wire_18;
	wire [3 : 0] fresh_wire_19;
	wire [0 : 0] fresh_wire_20;
	wire [0 : 0] fresh_wire_21;
	wire [0 : 0] fresh_wire_22;
	wire [0 : 0] fresh_wire_23;
	wire [0 : 0] fresh_wire_24;
	wire [0 : 0] fresh_wire_25;
	wire [0 : 0] fresh_wire_26;
	wire [0 : 0] fresh_wire_27;
	wire [0 : 0] fresh_wire_28;
	wire [0 : 0] fresh_wire_29;
	wire [0 : 0] fresh_wire_30;
	wire [0 : 0] fresh_wire_31;
	wire [0 : 0] fresh_wire_32;
	wire [0 : 0] fresh_wire_33;
	wire [0 : 0] fresh_wire_34;
	wire [0 : 0] fresh_wire_35;
	wire [0 : 0] fresh_wire_36;
	wire [0 : 0] fresh_wire_37;
	wire [0 : 0] fresh_wire_38;
	wire [0 : 0] fresh_wire_39;
	wire [0 : 0] fresh_wire_40;
	wire [0 : 0] fresh_wire_41;
	wire [0 : 0] fresh_wire_42;
	wire [0 : 0] fresh_wire_43;
	wire [0 : 0] fresh_wire_44;
	wire [0 : 0] fresh_wire_45;
	wire [0 : 0] fresh_wire_46;
	wire [0 : 0] fresh_wire_47;
	wire [0 : 0] fresh_wire_48;
	wire [0 : 0] fresh_wire_49;
	wire [0 : 0] fresh_wire_50;
	wire [0 : 0] fresh_wire_51;
	wire [0 : 0] fresh_wire_52;
	wire [0 : 0] fresh_wire_53;
	wire [0 : 0] fresh_wire_54;
	wire [0 : 0] fresh_wire_55;
	wire [0 : 0] fresh_wire_56;
	wire [0 : 0] fresh_wire_57;
	wire [0 : 0] fresh_wire_58;
	wire [0 : 0] fresh_wire_59;
	wire [0 : 0] fresh_wire_60;
	wire [0 : 0] fresh_wire_61;
	wire [0 : 0] fresh_wire_62;
	wire [0 : 0] fresh_wire_63;
	wire [0 : 0] fresh_wire_64;
	wire [0 : 0] fresh_wire_65;
	wire [0 : 0] fresh_wire_66;
	wire [0 : 0] fresh_wire_67;
	wire [0 : 0] fresh_wire_68;
	wire [0 : 0] fresh_wire_69;
	wire [0 : 0] fresh_wire_70;
	wire [0 : 0] fresh_wire_71;
	wire [0 : 0] fresh_wire_72;
	wire [0 : 0] fresh_wire_73;
	wire [0 : 0] fresh_wire_74;
	wire [0 : 0] fresh_wire_75;
	wire [0 : 0] fresh_wire_76;
	wire [0 : 0] fresh_wire_77;
	wire [0 : 0] fresh_wire_78;
	wire [0 : 0] fresh_wire_79;
	wire [0 : 0] fresh_wire_80;
	wire [0 : 0] fresh_wire_81;
	wire [0 : 0] fresh_wire_82;
	wire [0 : 0] fresh_wire_83;
	wire [0 : 0] fresh_wire_84;
	wire [0 : 0] fresh_wire_85;
	wire [0 : 0] fresh_wire_86;
	wire [0 : 0] fresh_wire_87;
	wire [0 : 0] fresh_wire_88;
	wire [0 : 0] fresh_wire_89;
	wire [0 : 0] fresh_wire_90;
	wire [0 : 0] fresh_wire_91;
	wire [0 : 0] fresh_wire_92;
	wire [0 : 0] fresh_wire_93;
	wire [0 : 0] fresh_wire_94;
	wire [0 : 0] fresh_wire_95;
	wire [0 : 0] fresh_wire_96;
	wire [0 : 0] fresh_wire_97;
	wire [0 : 0] fresh_wire_98;
	wire [0 : 0] fresh_wire_99;
	wire [0 : 0] fresh_wire_100;
	wire [0 : 0] fresh_wire_101;
	wire [0 : 0] fresh_wire_102;
	wire [0 : 0] fresh_wire_103;
	wire [0 : 0] fresh_wire_104;
	wire [0 : 0] fresh_wire_105;
	wire [0 : 0] fresh_wire_106;
	wire [0 : 0] fresh_wire_107;
	wire [0 : 0] fresh_wire_108;
	wire [0 : 0] fresh_wire_109;
	wire [0 : 0] fresh_wire_110;
	wire [0 : 0] fresh_wire_111;
	wire [0 : 0] fresh_wire_112;
	wire [0 : 0] fresh_wire_113;
	wire [0 : 0] fresh_wire_114;
	wire [0 : 0] fresh_wire_115;
	wire [0 : 0] fresh_wire_116;
	wire [0 : 0] fresh_wire_117;
	wire [0 : 0] fresh_wire_118;
	wire [0 : 0] fresh_wire_119;
	wire [0 : 0] fresh_wire_120;
	wire [0 : 0] fresh_wire_121;
	wire [0 : 0] fresh_wire_122;
	wire [0 : 0] fresh_wire_123;
	wire [0 : 0] fresh_wire_124;
	wire [0 : 0] fresh_wire_125;
	wire [0 : 0] fresh_wire_126;
	wire [0 : 0] fresh_wire_127;
	wire [0 : 0] fresh_wire_128;
	wire [0 : 0] fresh_wire_129;
	wire [0 : 0] fresh_wire_130;
	wire [0 : 0] fresh_wire_131;
	wire [0 : 0] fresh_wire_132;
	wire [0 : 0] fresh_wire_133;
	wire [0 : 0] fresh_wire_134;
	wire [0 : 0] fresh_wire_135;
	wire [0 : 0] fresh_wire_136;
	wire [0 : 0] fresh_wire_137;
	wire [0 : 0] fresh_wire_138;
	wire [0 : 0] fresh_wire_139;
	wire [0 : 0] fresh_wire_140;
	wire [0 : 0] fresh_wire_141;
	wire [0 : 0] fresh_wire_142;
	wire [0 : 0] fresh_wire_143;
	wire [0 : 0] fresh_wire_144;
	wire [0 : 0] fresh_wire_145;
	wire [0 : 0] fresh_wire_146;
	wire [0 : 0] fresh_wire_147;
	wire [0 : 0] fresh_wire_148;
	wire [0 : 0] fresh_wire_149;
	wire [0 : 0] fresh_wire_150;
	wire [0 : 0] fresh_wire_151;
	wire [0 : 0] fresh_wire_152;
	wire [0 : 0] fresh_wire_153;
	wire [12 : 0] fresh_wire_154;
	wire [16 : 0] fresh_wire_155;
	wire [33 : 0] fresh_wire_156;
	wire [33 : 0] fresh_wire_157;
	wire [33 : 0] fresh_wire_158;
	wire [33 : 0] fresh_wire_159;
	wire [0 : 0] fresh_wire_160;
	wire [0 : 0] fresh_wire_161;
	wire [33 : 0] fresh_wire_162;
	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) aux_div_pad_port_cell(.PORT_ID_IN(fresh_wire_0),
.PORT_ID_OUT(aux_div_pad));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) cell_261940_const_replacement(.PORT_ID_OUT(fresh_wire_161));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(34'h000000002),
.PARAM_WIDTH(32'h00000022)) cell_261945_const_replacement(.PORT_ID_OUT(fresh_wire_162));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) clk_ext_in_port_cell(.PORT_ID_IN(clk_ext_in),
.PORT_ID_OUT(fresh_wire_1));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) clk_in_port_cell(.PORT_ID_IN(clk_in),
.PORT_ID_OUT(fresh_wire_2));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000020),
.PARAM_PORT_TYPE(2'h0)) config_addr_in_port_cell(.PORT_ID_IN(config_addr_in),
.PORT_ID_OUT(fresh_wire_3));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000020),
.PARAM_PORT_TYPE(2'h0)) config_data_in_port_cell(.PORT_ID_IN(config_data_in),
.PORT_ID_OUT(fresh_wire_4));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) ext_cki_jm_port_cell(.PORT_ID_IN(ext_cki_jm),
.PORT_ID_OUT(fresh_wire_6));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) ext_cki_port_cell(.PORT_ID_IN(ext_cki),
.PORT_ID_OUT(fresh_wire_5));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) ext_ckib_jm_port_cell(.PORT_ID_IN(ext_ckib_jm),
.PORT_ID_OUT(fresh_wire_8));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) ext_ckib_port_cell(.PORT_ID_IN(ext_ckib),
.PORT_ID_OUT(fresh_wire_7));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) ext_frefn_jm_port_cell(.PORT_ID_IN(ext_frefn_jm),
.PORT_ID_OUT(fresh_wire_10));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) ext_frefn_port_cell(.PORT_ID_IN(ext_frefn),
.PORT_ID_OUT(fresh_wire_9));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) ext_frefp_jm_port_cell(.PORT_ID_IN(ext_frefp_jm),
.PORT_ID_OUT(fresh_wire_12));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) ext_frefp_port_cell(.PORT_ID_IN(ext_frefp),
.PORT_ID_OUT(fresh_wire_11));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) ffeed_pad_port_cell(.PORT_ID_IN(fresh_wire_13),
.PORT_ID_OUT(ffeed_pad));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) fout_div_pad_port_cell(.PORT_ID_IN(fresh_wire_14),
.PORT_ID_OUT(fout_div_pad));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) fref_off_pad_port_cell(.PORT_ID_IN(fresh_wire_15),
.PORT_ID_OUT(fref_off_pad));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) frefn_out_jm_port_cell(.PORT_ID_IN(fresh_wire_16),
.PORT_ID_OUT(frefn_out_jm));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) frefp_out_jm_port_cell(.PORT_ID_IN(fresh_wire_17),
.PORT_ID_OUT(frefp_out_jm));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h0000000d),
.PARAM_PORT_TYPE(2'h1)) lf_out_port_cell(.PORT_ID_IN(fresh_wire_18),
.PORT_ID_OUT(lf_out));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(13'h0000),
.PARAM_WIDTH(32'h0000000d)) mdll_top$self_lf_out(.PORT_ID_OUT(fresh_wire_154));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000004),
.PARAM_PORT_TYPE(2'h1)) mdllout_pad_port_cell(.PORT_ID_IN(fresh_wire_19),
.PORT_ID_OUT(mdllout_pad));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T0_in_port_cell(.PORT_ID_IN(pad_S0_T0_in),
.PORT_ID_OUT(fresh_wire_20));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T0_out_port_cell(.PORT_ID_IN(fresh_wire_21),
.PORT_ID_OUT(pad_S0_T0_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T10_in_port_cell(.PORT_ID_IN(pad_S0_T10_in),
.PORT_ID_OUT(fresh_wire_22));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T10_out_port_cell(.PORT_ID_IN(fresh_wire_23),
.PORT_ID_OUT(pad_S0_T10_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T11_in_port_cell(.PORT_ID_IN(pad_S0_T11_in),
.PORT_ID_OUT(fresh_wire_24));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T11_out_port_cell(.PORT_ID_IN(fresh_wire_25),
.PORT_ID_OUT(pad_S0_T11_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T12_in_port_cell(.PORT_ID_IN(pad_S0_T12_in),
.PORT_ID_OUT(fresh_wire_26));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T12_out_port_cell(.PORT_ID_IN(fresh_wire_27),
.PORT_ID_OUT(pad_S0_T12_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T13_in_port_cell(.PORT_ID_IN(pad_S0_T13_in),
.PORT_ID_OUT(fresh_wire_28));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T13_out_port_cell(.PORT_ID_IN(fresh_wire_29),
.PORT_ID_OUT(pad_S0_T13_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T14_in_port_cell(.PORT_ID_IN(pad_S0_T14_in),
.PORT_ID_OUT(fresh_wire_30));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T14_out_port_cell(.PORT_ID_IN(fresh_wire_31),
.PORT_ID_OUT(pad_S0_T14_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T15_in_port_cell(.PORT_ID_IN(pad_S0_T15_in),
.PORT_ID_OUT(fresh_wire_32));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T15_out_port_cell(.PORT_ID_IN(fresh_wire_33),
.PORT_ID_OUT(pad_S0_T15_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T1_in_port_cell(.PORT_ID_IN(pad_S0_T1_in),
.PORT_ID_OUT(fresh_wire_34));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T1_out_port_cell(.PORT_ID_IN(fresh_wire_35),
.PORT_ID_OUT(pad_S0_T1_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T2_in_port_cell(.PORT_ID_IN(pad_S0_T2_in),
.PORT_ID_OUT(fresh_wire_36));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T2_out_port_cell(.PORT_ID_IN(fresh_wire_37),
.PORT_ID_OUT(pad_S0_T2_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T3_in_port_cell(.PORT_ID_IN(pad_S0_T3_in),
.PORT_ID_OUT(fresh_wire_38));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T3_out_port_cell(.PORT_ID_IN(fresh_wire_39),
.PORT_ID_OUT(pad_S0_T3_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T4_in_port_cell(.PORT_ID_IN(pad_S0_T4_in),
.PORT_ID_OUT(fresh_wire_40));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T4_out_port_cell(.PORT_ID_IN(fresh_wire_41),
.PORT_ID_OUT(pad_S0_T4_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T5_in_port_cell(.PORT_ID_IN(pad_S0_T5_in),
.PORT_ID_OUT(fresh_wire_42));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T5_out_port_cell(.PORT_ID_IN(fresh_wire_43),
.PORT_ID_OUT(pad_S0_T5_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T6_in_port_cell(.PORT_ID_IN(pad_S0_T6_in),
.PORT_ID_OUT(fresh_wire_44));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T6_out_port_cell(.PORT_ID_IN(fresh_wire_45),
.PORT_ID_OUT(pad_S0_T6_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T7_in_port_cell(.PORT_ID_IN(pad_S0_T7_in),
.PORT_ID_OUT(fresh_wire_46));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T7_out_port_cell(.PORT_ID_IN(fresh_wire_47),
.PORT_ID_OUT(pad_S0_T7_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T8_in_port_cell(.PORT_ID_IN(pad_S0_T8_in),
.PORT_ID_OUT(fresh_wire_48));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T8_out_port_cell(.PORT_ID_IN(fresh_wire_49),
.PORT_ID_OUT(pad_S0_T8_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S0_T9_in_port_cell(.PORT_ID_IN(pad_S0_T9_in),
.PORT_ID_OUT(fresh_wire_50));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S0_T9_out_port_cell(.PORT_ID_IN(fresh_wire_51),
.PORT_ID_OUT(pad_S0_T9_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T0_in_port_cell(.PORT_ID_IN(pad_S1_T0_in),
.PORT_ID_OUT(fresh_wire_52));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T0_out_port_cell(.PORT_ID_IN(fresh_wire_53),
.PORT_ID_OUT(pad_S1_T0_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T10_in_port_cell(.PORT_ID_IN(pad_S1_T10_in),
.PORT_ID_OUT(fresh_wire_54));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T10_out_port_cell(.PORT_ID_IN(fresh_wire_55),
.PORT_ID_OUT(pad_S1_T10_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T11_in_port_cell(.PORT_ID_IN(pad_S1_T11_in),
.PORT_ID_OUT(fresh_wire_56));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T11_out_port_cell(.PORT_ID_IN(fresh_wire_57),
.PORT_ID_OUT(pad_S1_T11_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T12_in_port_cell(.PORT_ID_IN(pad_S1_T12_in),
.PORT_ID_OUT(fresh_wire_58));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T12_out_port_cell(.PORT_ID_IN(fresh_wire_59),
.PORT_ID_OUT(pad_S1_T12_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T13_in_port_cell(.PORT_ID_IN(pad_S1_T13_in),
.PORT_ID_OUT(fresh_wire_60));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T13_out_port_cell(.PORT_ID_IN(fresh_wire_61),
.PORT_ID_OUT(pad_S1_T13_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T14_in_port_cell(.PORT_ID_IN(pad_S1_T14_in),
.PORT_ID_OUT(fresh_wire_62));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T14_out_port_cell(.PORT_ID_IN(fresh_wire_63),
.PORT_ID_OUT(pad_S1_T14_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T15_in_port_cell(.PORT_ID_IN(pad_S1_T15_in),
.PORT_ID_OUT(fresh_wire_64));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T15_out_port_cell(.PORT_ID_IN(fresh_wire_65),
.PORT_ID_OUT(pad_S1_T15_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T1_in_port_cell(.PORT_ID_IN(pad_S1_T1_in),
.PORT_ID_OUT(fresh_wire_66));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T1_out_port_cell(.PORT_ID_IN(fresh_wire_67),
.PORT_ID_OUT(pad_S1_T1_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T2_in_port_cell(.PORT_ID_IN(pad_S1_T2_in),
.PORT_ID_OUT(fresh_wire_68));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T2_out_port_cell(.PORT_ID_IN(fresh_wire_69),
.PORT_ID_OUT(pad_S1_T2_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T3_in_port_cell(.PORT_ID_IN(pad_S1_T3_in),
.PORT_ID_OUT(fresh_wire_70));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T3_out_port_cell(.PORT_ID_IN(fresh_wire_71),
.PORT_ID_OUT(pad_S1_T3_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T4_in_port_cell(.PORT_ID_IN(pad_S1_T4_in),
.PORT_ID_OUT(fresh_wire_72));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T4_out_port_cell(.PORT_ID_IN(fresh_wire_73),
.PORT_ID_OUT(pad_S1_T4_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T5_in_port_cell(.PORT_ID_IN(pad_S1_T5_in),
.PORT_ID_OUT(fresh_wire_74));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T5_out_port_cell(.PORT_ID_IN(fresh_wire_75),
.PORT_ID_OUT(pad_S1_T5_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T6_in_port_cell(.PORT_ID_IN(pad_S1_T6_in),
.PORT_ID_OUT(fresh_wire_76));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T6_out_port_cell(.PORT_ID_IN(fresh_wire_77),
.PORT_ID_OUT(pad_S1_T6_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T7_in_port_cell(.PORT_ID_IN(pad_S1_T7_in),
.PORT_ID_OUT(fresh_wire_78));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T7_out_port_cell(.PORT_ID_IN(fresh_wire_79),
.PORT_ID_OUT(pad_S1_T7_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T8_in_port_cell(.PORT_ID_IN(pad_S1_T8_in),
.PORT_ID_OUT(fresh_wire_80));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T8_out_port_cell(.PORT_ID_IN(fresh_wire_81),
.PORT_ID_OUT(pad_S1_T8_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S1_T9_in_port_cell(.PORT_ID_IN(pad_S1_T9_in),
.PORT_ID_OUT(fresh_wire_82));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S1_T9_out_port_cell(.PORT_ID_IN(fresh_wire_83),
.PORT_ID_OUT(pad_S1_T9_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T0_in_port_cell(.PORT_ID_IN(pad_S2_T0_in),
.PORT_ID_OUT(fresh_wire_84));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T0_out_port_cell(.PORT_ID_IN(fresh_wire_85),
.PORT_ID_OUT(pad_S2_T0_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T10_in_port_cell(.PORT_ID_IN(pad_S2_T10_in),
.PORT_ID_OUT(fresh_wire_86));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T10_out_port_cell(.PORT_ID_IN(fresh_wire_87),
.PORT_ID_OUT(pad_S2_T10_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T11_in_port_cell(.PORT_ID_IN(pad_S2_T11_in),
.PORT_ID_OUT(fresh_wire_88));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T11_out_port_cell(.PORT_ID_IN(fresh_wire_89),
.PORT_ID_OUT(pad_S2_T11_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T12_in_port_cell(.PORT_ID_IN(pad_S2_T12_in),
.PORT_ID_OUT(fresh_wire_90));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T12_out_port_cell(.PORT_ID_IN(fresh_wire_91),
.PORT_ID_OUT(pad_S2_T12_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T13_in_port_cell(.PORT_ID_IN(pad_S2_T13_in),
.PORT_ID_OUT(fresh_wire_92));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T13_out_port_cell(.PORT_ID_IN(fresh_wire_93),
.PORT_ID_OUT(pad_S2_T13_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T14_in_port_cell(.PORT_ID_IN(pad_S2_T14_in),
.PORT_ID_OUT(fresh_wire_94));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T14_out_port_cell(.PORT_ID_IN(fresh_wire_95),
.PORT_ID_OUT(pad_S2_T14_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T15_in_port_cell(.PORT_ID_IN(pad_S2_T15_in),
.PORT_ID_OUT(fresh_wire_96));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T15_out_port_cell(.PORT_ID_IN(fresh_wire_97),
.PORT_ID_OUT(pad_S2_T15_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T1_in_port_cell(.PORT_ID_IN(pad_S2_T1_in),
.PORT_ID_OUT(fresh_wire_98));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T1_out_port_cell(.PORT_ID_IN(fresh_wire_99),
.PORT_ID_OUT(pad_S2_T1_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T2_in_port_cell(.PORT_ID_IN(pad_S2_T2_in),
.PORT_ID_OUT(fresh_wire_100));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T2_out_port_cell(.PORT_ID_IN(fresh_wire_101),
.PORT_ID_OUT(pad_S2_T2_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T3_in_port_cell(.PORT_ID_IN(pad_S2_T3_in),
.PORT_ID_OUT(fresh_wire_102));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T3_out_port_cell(.PORT_ID_IN(fresh_wire_103),
.PORT_ID_OUT(pad_S2_T3_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T4_in_port_cell(.PORT_ID_IN(pad_S2_T4_in),
.PORT_ID_OUT(fresh_wire_104));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T4_out_port_cell(.PORT_ID_IN(fresh_wire_105),
.PORT_ID_OUT(pad_S2_T4_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T5_in_port_cell(.PORT_ID_IN(pad_S2_T5_in),
.PORT_ID_OUT(fresh_wire_106));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T5_out_port_cell(.PORT_ID_IN(fresh_wire_107),
.PORT_ID_OUT(pad_S2_T5_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T6_in_port_cell(.PORT_ID_IN(pad_S2_T6_in),
.PORT_ID_OUT(fresh_wire_108));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T6_out_port_cell(.PORT_ID_IN(fresh_wire_109),
.PORT_ID_OUT(pad_S2_T6_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T7_in_port_cell(.PORT_ID_IN(pad_S2_T7_in),
.PORT_ID_OUT(fresh_wire_110));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T7_out_port_cell(.PORT_ID_IN(fresh_wire_111),
.PORT_ID_OUT(pad_S2_T7_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T8_in_port_cell(.PORT_ID_IN(pad_S2_T8_in),
.PORT_ID_OUT(fresh_wire_112));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T8_out_port_cell(.PORT_ID_IN(fresh_wire_113),
.PORT_ID_OUT(pad_S2_T8_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S2_T9_in_port_cell(.PORT_ID_IN(pad_S2_T9_in),
.PORT_ID_OUT(fresh_wire_114));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S2_T9_out_port_cell(.PORT_ID_IN(fresh_wire_115),
.PORT_ID_OUT(pad_S2_T9_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T0_in_port_cell(.PORT_ID_IN(pad_S3_T0_in),
.PORT_ID_OUT(fresh_wire_116));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T0_out_port_cell(.PORT_ID_IN(fresh_wire_117),
.PORT_ID_OUT(pad_S3_T0_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T10_in_port_cell(.PORT_ID_IN(pad_S3_T10_in),
.PORT_ID_OUT(fresh_wire_118));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T10_out_port_cell(.PORT_ID_IN(fresh_wire_119),
.PORT_ID_OUT(pad_S3_T10_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T11_in_port_cell(.PORT_ID_IN(pad_S3_T11_in),
.PORT_ID_OUT(fresh_wire_120));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T11_out_port_cell(.PORT_ID_IN(fresh_wire_121),
.PORT_ID_OUT(pad_S3_T11_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T12_in_port_cell(.PORT_ID_IN(pad_S3_T12_in),
.PORT_ID_OUT(fresh_wire_122));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T12_out_port_cell(.PORT_ID_IN(fresh_wire_123),
.PORT_ID_OUT(pad_S3_T12_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T13_in_port_cell(.PORT_ID_IN(pad_S3_T13_in),
.PORT_ID_OUT(fresh_wire_124));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T13_out_port_cell(.PORT_ID_IN(fresh_wire_125),
.PORT_ID_OUT(pad_S3_T13_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T14_in_port_cell(.PORT_ID_IN(pad_S3_T14_in),
.PORT_ID_OUT(fresh_wire_126));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T14_out_port_cell(.PORT_ID_IN(fresh_wire_127),
.PORT_ID_OUT(pad_S3_T14_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T15_in_port_cell(.PORT_ID_IN(pad_S3_T15_in),
.PORT_ID_OUT(fresh_wire_128));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T15_out_port_cell(.PORT_ID_IN(fresh_wire_129),
.PORT_ID_OUT(pad_S3_T15_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T1_in_port_cell(.PORT_ID_IN(pad_S3_T1_in),
.PORT_ID_OUT(fresh_wire_130));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T1_out_port_cell(.PORT_ID_IN(fresh_wire_131),
.PORT_ID_OUT(pad_S3_T1_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T2_in_port_cell(.PORT_ID_IN(pad_S3_T2_in),
.PORT_ID_OUT(fresh_wire_132));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T2_out_port_cell(.PORT_ID_IN(fresh_wire_133),
.PORT_ID_OUT(pad_S3_T2_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T3_in_port_cell(.PORT_ID_IN(pad_S3_T3_in),
.PORT_ID_OUT(fresh_wire_134));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T3_out_port_cell(.PORT_ID_IN(fresh_wire_135),
.PORT_ID_OUT(pad_S3_T3_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T4_in_port_cell(.PORT_ID_IN(pad_S3_T4_in),
.PORT_ID_OUT(fresh_wire_136));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T4_out_port_cell(.PORT_ID_IN(fresh_wire_137),
.PORT_ID_OUT(pad_S3_T4_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T5_in_port_cell(.PORT_ID_IN(pad_S3_T5_in),
.PORT_ID_OUT(fresh_wire_138));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T5_out_port_cell(.PORT_ID_IN(fresh_wire_139),
.PORT_ID_OUT(pad_S3_T5_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T6_in_port_cell(.PORT_ID_IN(pad_S3_T6_in),
.PORT_ID_OUT(fresh_wire_140));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T6_out_port_cell(.PORT_ID_IN(fresh_wire_141),
.PORT_ID_OUT(pad_S3_T6_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T7_in_port_cell(.PORT_ID_IN(pad_S3_T7_in),
.PORT_ID_OUT(fresh_wire_142));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T7_out_port_cell(.PORT_ID_IN(fresh_wire_143),
.PORT_ID_OUT(pad_S3_T7_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T8_in_port_cell(.PORT_ID_IN(pad_S3_T8_in),
.PORT_ID_OUT(fresh_wire_144));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T8_out_port_cell(.PORT_ID_IN(fresh_wire_145),
.PORT_ID_OUT(pad_S3_T8_out));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) pad_S3_T9_in_port_cell(.PORT_ID_IN(pad_S3_T9_in),
.PORT_ID_OUT(fresh_wire_146));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) pad_S3_T9_out_port_cell(.PORT_ID_IN(fresh_wire_147),
.PORT_ID_OUT(pad_S3_T9_out));

	CELL_TYPE_ZEXT #(.PARAM_IN_WIDTH(32'h00000011),
.PARAM_OUT_WIDTH(32'h00000022)) pe_0x15$test_pe$test_pe_comp$test_mult_add$__DOLLAR__mul__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__1503$extendA(.PORT_ID_IN(fresh_wire_155),
.PORT_ID_OUT(fresh_wire_156));

	CELL_TYPE_MUL #(.PARAM_WIDTH(32'h00000022)) pe_0x15$test_pe$test_pe_comp$test_mult_add$__DOLLAR__mul__DOLLAR____FORWARD_SLASH__Users__FORWARD_SLASH__dillon__FORWARD_SLASH__CoreIRWorkspace__FORWARD_SLASH__CGRA_coreir__FORWARD_SLASH__cgra_with_config_ports__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__1503$op0(.PORT_ID_IN0(fresh_wire_157),
.PORT_ID_IN1(fresh_wire_158),
.PORT_ID_OUT(fresh_wire_159));

	CELL_TYPE_CONST #(.PARAM_INIT_VALUE(1'h0),
.PARAM_WIDTH(32'h00000001)) pe_0xFF__DOT__tile_id__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(.PORT_ID_OUT(fresh_wire_160));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) reset_in_port_cell(.PORT_ID_IN(reset_in),
.PORT_ID_OUT(fresh_wire_148));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) tck_port_cell(.PORT_ID_IN(tck),
.PORT_ID_OUT(fresh_wire_149));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) tdi_port_cell(.PORT_ID_IN(tdi),
.PORT_ID_OUT(fresh_wire_150));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h1)) tdo_port_cell(.PORT_ID_IN(fresh_wire_151),
.PORT_ID_OUT(tdo));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) tms_port_cell(.PORT_ID_IN(tms),
.PORT_ID_OUT(fresh_wire_152));

	CELL_TYPE_PORT #(.PARAM_OUT_WIDTH(32'h00000001),
.PARAM_PORT_TYPE(2'h0)) trst_n_port_cell(.PORT_ID_IN(trst_n),
.PORT_ID_OUT(fresh_wire_153));

	assign fresh_wire_0[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_13[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_14[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_15[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_16[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_17[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_18[ 0 ] = fresh_wire_154[ 0 ];
	assign fresh_wire_18[ 1 ] = fresh_wire_154[ 1 ];
	assign fresh_wire_18[ 2 ] = fresh_wire_154[ 2 ];
	assign fresh_wire_18[ 3 ] = fresh_wire_154[ 3 ];
	assign fresh_wire_18[ 4 ] = fresh_wire_154[ 4 ];
	assign fresh_wire_18[ 5 ] = fresh_wire_154[ 5 ];
	assign fresh_wire_18[ 6 ] = fresh_wire_154[ 6 ];
	assign fresh_wire_18[ 7 ] = fresh_wire_154[ 7 ];
	assign fresh_wire_18[ 8 ] = fresh_wire_154[ 8 ];
	assign fresh_wire_18[ 9 ] = fresh_wire_154[ 9 ];
	assign fresh_wire_18[ 10 ] = fresh_wire_154[ 10 ];
	assign fresh_wire_18[ 11 ] = fresh_wire_154[ 11 ];
	assign fresh_wire_18[ 12 ] = fresh_wire_154[ 12 ];
	assign fresh_wire_19[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_19[ 1 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_19[ 2 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_19[ 3 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_21[ 0 ] = fresh_wire_159[ 15 ];
	assign fresh_wire_23[ 0 ] = fresh_wire_159[ 5 ];
	assign fresh_wire_25[ 0 ] = fresh_wire_159[ 4 ];
	assign fresh_wire_27[ 0 ] = fresh_wire_159[ 3 ];
	assign fresh_wire_29[ 0 ] = fresh_wire_159[ 2 ];
	assign fresh_wire_31[ 0 ] = fresh_wire_159[ 1 ];
	assign fresh_wire_33[ 0 ] = fresh_wire_159[ 0 ];
	assign fresh_wire_35[ 0 ] = fresh_wire_159[ 14 ];
	assign fresh_wire_37[ 0 ] = fresh_wire_159[ 13 ];
	assign fresh_wire_39[ 0 ] = fresh_wire_159[ 12 ];
	assign fresh_wire_41[ 0 ] = fresh_wire_159[ 11 ];
	assign fresh_wire_43[ 0 ] = fresh_wire_159[ 10 ];
	assign fresh_wire_45[ 0 ] = fresh_wire_159[ 9 ];
	assign fresh_wire_47[ 0 ] = fresh_wire_159[ 8 ];
	assign fresh_wire_49[ 0 ] = fresh_wire_159[ 7 ];
	assign fresh_wire_51[ 0 ] = fresh_wire_159[ 6 ];
	assign fresh_wire_53[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_55[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_57[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_59[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_61[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_63[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_65[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_67[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_69[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_71[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_73[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_75[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_77[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_79[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_81[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_83[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_85[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_87[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_89[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_91[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_93[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_95[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_97[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_99[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_101[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_103[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_105[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_107[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_109[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_111[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_113[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_115[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_117[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_119[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_121[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_123[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_125[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_127[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_129[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_131[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_133[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_135[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_137[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_139[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_141[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_143[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_145[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_147[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_151[ 0 ] = fresh_wire_160[ 0 ];
	assign fresh_wire_155[ 0 ] = fresh_wire_96[ 0 ];
	assign fresh_wire_155[ 1 ] = fresh_wire_94[ 0 ];
	assign fresh_wire_155[ 2 ] = fresh_wire_92[ 0 ];
	assign fresh_wire_155[ 3 ] = fresh_wire_90[ 0 ];
	assign fresh_wire_155[ 4 ] = fresh_wire_88[ 0 ];
	assign fresh_wire_155[ 5 ] = fresh_wire_86[ 0 ];
	assign fresh_wire_155[ 6 ] = fresh_wire_114[ 0 ];
	assign fresh_wire_155[ 7 ] = fresh_wire_112[ 0 ];
	assign fresh_wire_155[ 8 ] = fresh_wire_110[ 0 ];
	assign fresh_wire_155[ 9 ] = fresh_wire_108[ 0 ];
	assign fresh_wire_155[ 10 ] = fresh_wire_106[ 0 ];
	assign fresh_wire_155[ 11 ] = fresh_wire_104[ 0 ];
	assign fresh_wire_155[ 12 ] = fresh_wire_102[ 0 ];
	assign fresh_wire_155[ 13 ] = fresh_wire_100[ 0 ];
	assign fresh_wire_155[ 14 ] = fresh_wire_98[ 0 ];
	assign fresh_wire_155[ 15 ] = fresh_wire_84[ 0 ];
	assign fresh_wire_155[ 16 ] = fresh_wire_161[ 0 ];
	assign fresh_wire_157[ 0 ] = fresh_wire_156[ 0 ];
	assign fresh_wire_157[ 1 ] = fresh_wire_156[ 1 ];
	assign fresh_wire_157[ 2 ] = fresh_wire_156[ 2 ];
	assign fresh_wire_157[ 3 ] = fresh_wire_156[ 3 ];
	assign fresh_wire_157[ 4 ] = fresh_wire_156[ 4 ];
	assign fresh_wire_157[ 5 ] = fresh_wire_156[ 5 ];
	assign fresh_wire_157[ 6 ] = fresh_wire_156[ 6 ];
	assign fresh_wire_157[ 7 ] = fresh_wire_156[ 7 ];
	assign fresh_wire_157[ 8 ] = fresh_wire_156[ 8 ];
	assign fresh_wire_157[ 9 ] = fresh_wire_156[ 9 ];
	assign fresh_wire_157[ 10 ] = fresh_wire_156[ 10 ];
	assign fresh_wire_157[ 11 ] = fresh_wire_156[ 11 ];
	assign fresh_wire_157[ 12 ] = fresh_wire_156[ 12 ];
	assign fresh_wire_157[ 13 ] = fresh_wire_156[ 13 ];
	assign fresh_wire_157[ 14 ] = fresh_wire_156[ 14 ];
	assign fresh_wire_157[ 15 ] = fresh_wire_156[ 15 ];
	assign fresh_wire_157[ 16 ] = fresh_wire_156[ 16 ];
	assign fresh_wire_157[ 17 ] = fresh_wire_156[ 17 ];
	assign fresh_wire_157[ 18 ] = fresh_wire_156[ 18 ];
	assign fresh_wire_157[ 19 ] = fresh_wire_156[ 19 ];
	assign fresh_wire_157[ 20 ] = fresh_wire_156[ 20 ];
	assign fresh_wire_157[ 21 ] = fresh_wire_156[ 21 ];
	assign fresh_wire_157[ 22 ] = fresh_wire_156[ 22 ];
	assign fresh_wire_157[ 23 ] = fresh_wire_156[ 23 ];
	assign fresh_wire_157[ 24 ] = fresh_wire_156[ 24 ];
	assign fresh_wire_157[ 25 ] = fresh_wire_156[ 25 ];
	assign fresh_wire_157[ 26 ] = fresh_wire_156[ 26 ];
	assign fresh_wire_157[ 27 ] = fresh_wire_156[ 27 ];
	assign fresh_wire_157[ 28 ] = fresh_wire_156[ 28 ];
	assign fresh_wire_157[ 29 ] = fresh_wire_156[ 29 ];
	assign fresh_wire_157[ 30 ] = fresh_wire_156[ 30 ];
	assign fresh_wire_157[ 31 ] = fresh_wire_156[ 31 ];
	assign fresh_wire_157[ 32 ] = fresh_wire_156[ 32 ];
	assign fresh_wire_157[ 33 ] = fresh_wire_156[ 33 ];
	assign fresh_wire_158[ 0 ] = fresh_wire_162[ 0 ];
	assign fresh_wire_158[ 1 ] = fresh_wire_162[ 1 ];
	assign fresh_wire_158[ 2 ] = fresh_wire_162[ 2 ];
	assign fresh_wire_158[ 3 ] = fresh_wire_162[ 3 ];
	assign fresh_wire_158[ 4 ] = fresh_wire_162[ 4 ];
	assign fresh_wire_158[ 5 ] = fresh_wire_162[ 5 ];
	assign fresh_wire_158[ 6 ] = fresh_wire_162[ 6 ];
	assign fresh_wire_158[ 7 ] = fresh_wire_162[ 7 ];
	assign fresh_wire_158[ 8 ] = fresh_wire_162[ 8 ];
	assign fresh_wire_158[ 9 ] = fresh_wire_162[ 9 ];
	assign fresh_wire_158[ 10 ] = fresh_wire_162[ 10 ];
	assign fresh_wire_158[ 11 ] = fresh_wire_162[ 11 ];
	assign fresh_wire_158[ 12 ] = fresh_wire_162[ 12 ];
	assign fresh_wire_158[ 13 ] = fresh_wire_162[ 13 ];
	assign fresh_wire_158[ 14 ] = fresh_wire_162[ 14 ];
	assign fresh_wire_158[ 15 ] = fresh_wire_162[ 15 ];
	assign fresh_wire_158[ 16 ] = fresh_wire_162[ 16 ];
	assign fresh_wire_158[ 17 ] = fresh_wire_162[ 17 ];
	assign fresh_wire_158[ 18 ] = fresh_wire_162[ 18 ];
	assign fresh_wire_158[ 19 ] = fresh_wire_162[ 19 ];
	assign fresh_wire_158[ 20 ] = fresh_wire_162[ 20 ];
	assign fresh_wire_158[ 21 ] = fresh_wire_162[ 21 ];
	assign fresh_wire_158[ 22 ] = fresh_wire_162[ 22 ];
	assign fresh_wire_158[ 23 ] = fresh_wire_162[ 23 ];
	assign fresh_wire_158[ 24 ] = fresh_wire_162[ 24 ];
	assign fresh_wire_158[ 25 ] = fresh_wire_162[ 25 ];
	assign fresh_wire_158[ 26 ] = fresh_wire_162[ 26 ];
	assign fresh_wire_158[ 27 ] = fresh_wire_162[ 27 ];
	assign fresh_wire_158[ 28 ] = fresh_wire_162[ 28 ];
	assign fresh_wire_158[ 29 ] = fresh_wire_162[ 29 ];
	assign fresh_wire_158[ 30 ] = fresh_wire_162[ 30 ];
	assign fresh_wire_158[ 31 ] = fresh_wire_162[ 31 ];
	assign fresh_wire_158[ 32 ] = fresh_wire_162[ 32 ];
	assign fresh_wire_158[ 33 ] = fresh_wire_162[ 33 ];
endmodule

